module data_concat_tb #()
(

);


endmodule