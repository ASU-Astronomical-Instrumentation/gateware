`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 02/08/2021 02:10:06 PM
// Design Name: 
// Module Name: ddc_top
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module ddc_top #(
        //parameter BINS = 10;
    )
    (
    input wire clk, a_reset, s_axis_a_tvalid, s_axis_b_tvalid,
    input wire [31:0] x0_real_res1, x0_im_res1, x0_real_res2, x0_im_res2,
    input wire [31:0] x1_real_res1, x1_im_res1, x1_real_res2, x1_im_res2,
    input wire [31:0] x2_real_res1, x2_im_res1, x2_real_res2, x2_im_res2,
    input wire [31:0] x3_real_res1, x3_im_res1, x3_real_res2, x3_im_res2,
    output reg [79:0] x0_real_res1_out, x0_im_res1_out
    );
    
//----------------------------------------------
//------------ INTERANAL SIGNALS ---------------    
//----------------------------------------------
    reg [31:0] counter;
    wire [79:0] cmult_x0_real_res1, cmult_x0_im_res1, cmult_x0_real_res2, cmult_x0_im_res2;
    wire [79:0] cmult_x1_real_res1, cmult_x1_im_res1, cmult_x1_real_res2, cmult_x1_im_res2;
    wire [79:0] cmult_x2_real_res1, cmult_x2_im_res1, cmult_x2_real_res2, cmult_x2_im_res2;
    wire [79:0] cmult_x3_real_res1, cmult_x3_im_res1, cmult_x3_real_res2, cmult_x3_im_res2;

    
    //complex mult output valid signal
    wire dout_tvalid_x0_real_res1, dout_tvalid_x0_im_res1, dout_tvalid_x0_real_res2, dout_tvalid_x0_im_res2;
    wire dout_tvalid_x1_real_res1, dout_tvalid_x1_im_res1, dout_tvalid_x1_real_res2, dout_tvalid_x1_im_res2;
    wire dout_tvalid_x2_real_res1, dout_tvalid_x2_im_res1, dout_tvalid_x2_real_res2, dout_tvalid_x2_im_res2;
    wire dout_tvalid_x3_real_res1, dout_tvalid_x3_im_res1, dout_tvalid_x3_real_res2, dout_tvalid_x3_im_res2;

    //LUT values 
    reg [31:0] LUT_x0_real_res1, LUT_x0_im_res1, LUT_x0_real_res2, LUT_x0_im_res2;
    reg [31:0] LUT_x1_real_res1, LUT_x1_im_res1, LUT_x1_real_res2, LUT_x1_im_res2;
    reg [31:0] LUT_x2_real_res1, LUT_x2_im_res1, LUT_x2_real_res2, LUT_x2_im_res2;
    reg [31:0] LUT_x3_real_res1, LUT_x3_im_res1, LUT_x3_real_res2, LUT_x3_im_res2;
    reg aclken;
    
//----------------------------------------------
//--------- INTERANAL DELAY SIGNALS ------------    
//----------------------------------------------
    //LUT delays
    reg [31:0] LUT_x0_real_res1_d1, LUT_x0_im_res1_d1, LUT_x0_real_res2_d1, LUT_x0_im_res2_d1;
    reg [31:0] LUT_x1_real_res1_d1, LUT_x1_im_res1_d1, LUT_x1_real_res2_d1, LUT_x1_im_res2_d1;
    reg [31:0] LUT_x2_real_res1_d1, LUT_x2_im_res1_d1, LUT_x2_real_res2_d1, LUT_x2_im_res2_d1;
    reg [31:0] LUT_x3_real_res1_d1, LUT_x3_im_res1_d1, LUT_x3_real_res2_d1, LUT_x3_im_res2_d1;
    
    //input PFB delays
    reg [31:0] x0_real_res1_d1, x0_real_res1_d2, x0_im_res1_d1, x0_im_res1_d2;
    reg [31:0] x0_real_res2_d1, x0_real_res2_d2, x0_im_res2_d1, x0_im_res2_d2;
    reg [31:0] x1_real_res1_d1, x1_real_res1_d2, x1_im_res1_d1, x1_im_res1_d2;
    reg [31:0] x1_real_res2_d1, x1_real_res2_d2, x1_im_res2_d1, x1_im_res2_d2;
    reg [31:0] x2_real_res1_d1, x2_real_res1_d2, x2_im_res1_d1, x2_im_res1_d2;
    reg [31:0] x2_real_res2_d1, x2_real_res2_d2, x2_im_res2_d1, x2_im_res2_d2;
    reg [31:0] x3_real_res1_d1, x3_real_res1_d2, x3_im_res1_d1, x3_im_res1_d2;
    reg [31:0] x3_real_res2_d1, x3_real_res2_d2, x3_im_res2_d1, x3_im_res2_d2;    
        
//----------------------------------------------
//-------------- DATA HANDLING -----------------    
//----------------------------------------------
    
    always @ (posedge clk or negedge a_reset)
        if (a_reset) begin
            x0_real_res1_out <= 80'd0;
            x0_im_res1_out <= 80'd0;
        end
        else begin
            x0_real_res1_out <= cmult_x0_real_res1;
            x0_im_res1_out <= cmult_x0_im_res1;
        end
   
   //COUNTER 
   always @ (posedge clk or negedge a_reset) 
        if (~a_reset) begin
            counter <= 31'd0;
            aclken <= 1'b0;
        end
        else if (counter == 256) begin
            counter <= 31'd1;
            aclken <= 1'b0;
        end else begin
            counter <= counter + 1;
            aclken <= 1'b1;
        end
        
    //delay input signal from PFB for cmult    
    always @ (posedge clk or negedge a_reset)
        if (~a_reset) begin
            //x0, resonator 1
            x0_real_res1_d1 <= 0;
            x0_real_res1_d2 <= 0;
            x0_im_res1_d1 <= 0;
            x0_im_res1_d2 <= 0;
            //x0, resonator 2
            x0_real_res2_d1 <= 0;
            x0_real_res2_d2 <= 0;
            x0_im_res2_d1 <= 0;
            x0_im_res2_d2 <= 0;
            //x1, resonator 1
            x1_real_res1_d1 <= 0;
            x1_real_res1_d2 <= 0;
            x1_im_res1_d1 <= 0;
            x1_im_res1_d2 <= 0;
            //x1, resonator 2
            x1_real_res2_d1 <= 0;
            x1_real_res2_d2 <= 0;
            x1_im_res2_d1 <= 0;
            x1_im_res2_d2 <= 0;
            //x2, resonator 1
            x2_real_res1_d1 <= 0;
            x2_real_res1_d2 <= 0;
            x2_im_res1_d1 <= 0;
            x2_im_res1_d2 <= 0;
            //x2, resonator 2
            x2_real_res2_d1 <= 0;
            x2_real_res2_d2 <= 0;
            x2_im_res2_d1 <= 0;
            x2_im_res2_d2 <= 0;            
            //x3, resonator 1
            x3_real_res1_d1 <= 0;
            x3_real_res1_d2 <= 0;
            x3_im_res1_d1 <= 0;
            x3_im_res1_d2 <= 0;
            //x3, resonator 2
            x3_real_res2_d1 <= 0;
            x3_real_res2_d2 <= 0;
            x3_im_res2_d1 <= 0;
            x3_im_res2_d2 <= 0;
        end
        else begin
            //x0, resonator 1
            x0_real_res1_d1 <= x0_real_res1;
            x0_real_res1_d2 <= x0_real_res1_d1;
            x0_im_res1_d1 <= x0_im_res1;
            x0_im_res1_d2 <= x0_im_res1_d1;
            //x0, resonator 2
            x0_real_res2_d1 <= x0_real_res2;
            x0_real_res2_d2 <= x0_real_res2_d1;
            x0_im_res2_d1 <= x0_im_res2;
            x0_im_res2_d2 <= x0_im_res2_d1;
            //x1, resonator 1
            x1_real_res1_d1 <= x1_real_res1;
            x1_real_res1_d2 <= x1_real_res1_d1;
            x1_im_res1_d1 <= x1_im_res1;
            x1_im_res1_d2 <= x1_im_res1_d1;
            //x1, resonator 2
            x1_real_res2_d1 <= x1_real_res2;
            x1_real_res2_d2 <= x1_real_res2_d1;
            x1_im_res2_d1 <= x1_im_res2;
            x1_im_res2_d2 <= x1_im_res2_d1;
            //x2, resonator 1
            x2_real_res1_d1 <= x2_real_res1;
            x2_real_res1_d2 <= x2_real_res1_d1;
            x2_im_res1_d1 <= x2_im_res1;
            x2_im_res1_d2 <= x2_im_res1_d1;
            //x2, resonator 2
            x2_real_res2_d1 <= x2_real_res2;
            x2_real_res2_d2 <= x2_real_res2_d1;
            x2_im_res2_d1 <= x2_im_res2;
            x2_im_res2_d2 <= x2_im_res2_d1;
            //x3, resonator 1
            x3_real_res1_d1 <= x3_real_res1;
            x3_real_res1_d2 <= x3_real_res1_d1;
            x3_im_res1_d1 <= x3_im_res1;
            x3_im_res1_d2 <= x3_im_res1_d1;
            //x3, resonator 2
            x3_real_res2_d1 <= x3_real_res2;
            x3_real_res2_d2 <= x3_real_res2_d1;
            x3_im_res2_d1 <= x3_im_res2;
            x3_im_res2_d2 <= x3_im_res2_d1;
        end

//------------------------------------------------
//---------- COMPLEX MULTIPLICATION --------------
//------------------------------------------------   
    //x0 complex multiplies 
   cmpy_0 u_x0_real_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x0_real_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x0_real_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x0_real_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x0_real_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x0_im_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                            // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x0_im_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x0_im_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x0_im_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x0_im_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x0_real_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x0_real_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x0_real_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x0_real_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x0_real_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x0_im_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x0_im_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x0_im_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x0_im_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x0_im_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    //x1 complex multiplies 
       cmpy_0 u_x1_real_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x1_real_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x1_real_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x1_real_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x1_real_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x1_im_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                            // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x1_im_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x1_im_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x1_im_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x1_im_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x1_real_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x1_real_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x1_real_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x1_real_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x1_real_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x1_im_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x1_im_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x1_im_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x1_im_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x1_im_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    //x2 complex multiplies 
       cmpy_0 u_x2_real_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x2_real_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x2_real_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x2_real_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x2_real_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x2_im_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                            // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x2_im_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x2_im_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x2_im_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x2_im_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x2_real_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x2_real_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x2_real_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x2_real_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x2_real_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x2_im_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x2_im_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x2_im_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x2_im_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x2_im_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    //x3 complex multiplies 
       cmpy_0 u_x3_real_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x3_real_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x3_real_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x3_real_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x3_real_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x3_im_res1 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                            // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x3_im_res1_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x3_im_res1_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x3_im_res1),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x3_im_res1)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x3_real_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x3_real_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x3_real_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x3_real_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x3_real_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );
    
    cmpy_0 u_x3_im_res2 (
        .aclk(clk),  
        .aclken(1'b1),                          // input wire aclken
        .aresetn(a_reset),                             // input wire aclk
        .s_axis_a_tvalid(s_axis_a_tvalid),        // input wire s_axis_a_tvalid
        .s_axis_a_tdata(x3_im_res2_d2),          // input wire [31 : 0] s_axis_a_tdata
        .s_axis_b_tvalid(s_axis_b_tvalid),        // input wire s_axis_b_tvalid
        .s_axis_b_tdata(LUT_x3_im_res2_d1),          // input wire [31 : 0] s_axis_b_tdata
        .m_axis_dout_tvalid(dout_tvalid_x3_im_res2),  // output wire m_axis_dout_tvalid
        .m_axis_dout_tdata(cmult_x3_im_res2)    // output wire [79 : 0] m_axis_dout_tdata
    );

//----------------------------------------------
//----------- DELAY LUT SIGNALS ----------------    
//----------------------------------------------
    always @ (posedge clk or negedge a_reset) 
        if (~a_reset) begin
            //x0
            LUT_x0_real_res1_d1 <= 0;
            LUT_x0_im_res1_d1 <= 0;
            LUT_x0_real_res2_d1 <= 0;
            LUT_x0_im_res2_d1 <= 0;
            //x1
            LUT_x1_real_res1_d1 <= 0;
            LUT_x1_im_res1_d1 <= 0;
            LUT_x1_real_res2_d1 <= 0;
            LUT_x1_im_res2_d1 <= 0;
            //x2
            LUT_x2_real_res1_d1 <= 0;
            LUT_x2_im_res1_d1 <= 0;
            LUT_x2_real_res2_d1 <= 0;
            LUT_x2_im_res2_d1 <= 0;
            //x3
            LUT_x3_real_res1_d1 <= 0;
            LUT_x3_im_res1_d1 <= 0;
            LUT_x3_real_res2_d1 <= 0;
            LUT_x3_im_res2_d1 <= 0;
        end
        else begin
            //x0
            LUT_x0_real_res1_d1 <= LUT_x0_real_res1;
            LUT_x0_im_res1_d1 <= LUT_x0_im_res1;
            LUT_x0_real_res2_d1 <= LUT_x0_real_res2;
            LUT_x0_im_res2_d1 <= LUT_x0_im_res2;
            //x1
            LUT_x1_real_res1_d1 <= LUT_x1_real_res1;
            LUT_x1_im_res1_d1 <= LUT_x1_im_res1;
            LUT_x1_real_res2_d1 <= LUT_x1_real_res2;
            LUT_x1_im_res2_d1 <= LUT_x1_im_res2;
            //x2
            LUT_x2_real_res1_d1 <= LUT_x2_real_res1;
            LUT_x2_im_res1_d1 <= LUT_x2_im_res1;
            LUT_x2_real_res2_d1 <= LUT_x2_real_res2;
            LUT_x2_im_res2_d1 <= LUT_x2_im_res2;
            //x3
            LUT_x3_real_res1_d1 <= LUT_x3_real_res1;
            LUT_x3_im_res1_d1 <= LUT_x3_im_res1;
            LUT_x3_real_res2_d1 <= LUT_x3_real_res2;
            LUT_x3_im_res2_d1 <= LUT_x3_im_res2;
        end
        
//---------------------------------------------------
//------------ LUT INSTANTIATION --------------------
//---------------------------------------------------        
    
    //X0, resonator 1, real    
    always @(*) begin
        case(counter) 
            'd1: LUT_x0_real_res1 = 1;
            'd2: LUT_x0_real_res1 = 2;
            'd3: LUT_x0_real_res1 = 3;
            'd4: LUT_x0_real_res1 = 4;
            'd5: LUT_x0_real_res1 = 5;
            'd6: LUT_x0_real_res1 = 6;
            'd7: LUT_x0_real_res1 = 7;
            'd8: LUT_x0_real_res1 = 8;
            'd9: LUT_x0_real_res1 = 9;
            'd10: LUT_x0_real_res1 = 10;
            'd11: LUT_x0_real_res1 = 11;
            'd12: LUT_x0_real_res1 = 12;
            'd13: LUT_x0_real_res1 = 13;
            'd14: LUT_x0_real_res1 = 14;
            'd15: LUT_x0_real_res1 = 15;
            'd16: LUT_x0_real_res1 = 16;
            'd17: LUT_x0_real_res1 = 17;
            'd18: LUT_x0_real_res1 = 18;
            'd19: LUT_x0_real_res1 = 19;
            'd20: LUT_x0_real_res1 = 20;
            'd21: LUT_x0_real_res1 = 21;
            'd22: LUT_x0_real_res1 = 22;
            'd23: LUT_x0_real_res1 = 23;
            'd24: LUT_x0_real_res1 = 24;
            'd25: LUT_x0_real_res1 = 25;
            'd26: LUT_x0_real_res1 = 26;
            'd27: LUT_x0_real_res1 = 27;
            'd28: LUT_x0_real_res1 = 28;
            'd29: LUT_x0_real_res1 = 29;
            'd30: LUT_x0_real_res1 = 30;
            'd31: LUT_x0_real_res1 = 31;
            'd32: LUT_x0_real_res1 = 32;
            'd33: LUT_x0_real_res1 = 33;
            'd34: LUT_x0_real_res1 = 34;
            'd35: LUT_x0_real_res1 = 35;
            'd36: LUT_x0_real_res1 = 36;
            'd37: LUT_x0_real_res1 = 37;
            'd38: LUT_x0_real_res1 = 38;
            'd39: LUT_x0_real_res1 = 39;
            'd40: LUT_x0_real_res1 = 40;
            'd41: LUT_x0_real_res1 = 41;
            'd42: LUT_x0_real_res1 = 42;
            'd43: LUT_x0_real_res1 = 43;
            'd44: LUT_x0_real_res1 = 44;
            'd45: LUT_x0_real_res1 = 45;
            'd46: LUT_x0_real_res1 = 46;
            'd47: LUT_x0_real_res1 = 47;
            'd48: LUT_x0_real_res1 = 48;
            'd49: LUT_x0_real_res1 = 49;
            'd50: LUT_x0_real_res1 = 50;
            'd51: LUT_x0_real_res1 = 51;
            'd52: LUT_x0_real_res1 = 52;
            'd53: LUT_x0_real_res1 = 53;
            'd54: LUT_x0_real_res1 = 54;
            'd55: LUT_x0_real_res1 = 55;
            'd56: LUT_x0_real_res1 = 56;
            'd57: LUT_x0_real_res1 = 57;
            'd58: LUT_x0_real_res1 = 58;
            'd59: LUT_x0_real_res1 = 59;
            'd60: LUT_x0_real_res1 = 60;
            'd61: LUT_x0_real_res1 = 61;
            'd62: LUT_x0_real_res1 = 62;
            'd63: LUT_x0_real_res1 = 63;
            'd64: LUT_x0_real_res1 = 64;
            'd65: LUT_x0_real_res1 = 65;
            'd66: LUT_x0_real_res1 = 66;
            'd67: LUT_x0_real_res1 = 67;
            'd68: LUT_x0_real_res1 = 68;
            'd69: LUT_x0_real_res1 = 69;
            'd70: LUT_x0_real_res1 = 70;
            'd71: LUT_x0_real_res1 = 71;
            'd72: LUT_x0_real_res1 = 72;
            'd73: LUT_x0_real_res1 = 73;
            'd74: LUT_x0_real_res1 = 74;
            'd75: LUT_x0_real_res1 = 75;
            'd76: LUT_x0_real_res1 = 76;
            'd77: LUT_x0_real_res1 = 77;
            'd78: LUT_x0_real_res1 = 78;
            'd79: LUT_x0_real_res1 = 79;
            'd80: LUT_x0_real_res1 = 80;
            'd81: LUT_x0_real_res1 = 81;
            'd82: LUT_x0_real_res1 = 82;
            'd83: LUT_x0_real_res1 = 83;
            'd84: LUT_x0_real_res1 = 84;
            'd85: LUT_x0_real_res1 = 85;
            'd86: LUT_x0_real_res1 = 86;
            'd87: LUT_x0_real_res1 = 87;
            'd88: LUT_x0_real_res1 = 88;
            'd89: LUT_x0_real_res1 = 89;
            'd90: LUT_x0_real_res1 = 90;
            'd91: LUT_x0_real_res1 = 91;
            'd92: LUT_x0_real_res1 = 92;
            'd93: LUT_x0_real_res1 = 93;
            'd94: LUT_x0_real_res1 = 94;
            'd95: LUT_x0_real_res1 = 95;
            'd96: LUT_x0_real_res1 = 96;
            'd97: LUT_x0_real_res1 = 97;
            'd98: LUT_x0_real_res1 = 98;
            'd99: LUT_x0_real_res1 = 99;
            'd100: LUT_x0_real_res1 = 100;
            'd101: LUT_x0_real_res1 = 101;
            'd102: LUT_x0_real_res1 = 102;
            'd103: LUT_x0_real_res1 = 103;
            'd104: LUT_x0_real_res1 = 104;
            'd105: LUT_x0_real_res1 = 105;
            'd106: LUT_x0_real_res1 = 106;
            'd107: LUT_x0_real_res1 = 107;
            'd108: LUT_x0_real_res1 = 108;
            'd109: LUT_x0_real_res1 = 109;
            'd110: LUT_x0_real_res1 = 110;
            'd111: LUT_x0_real_res1 = 111;
            'd112: LUT_x0_real_res1 = 112;
            'd113: LUT_x0_real_res1 = 113;
            'd114: LUT_x0_real_res1 = 114;
            'd115: LUT_x0_real_res1 = 115;
            'd116: LUT_x0_real_res1 = 116;
            'd117: LUT_x0_real_res1 = 117;
            'd118: LUT_x0_real_res1 = 118;
            'd119: LUT_x0_real_res1 = 119;
            'd120: LUT_x0_real_res1 = 120;
            'd121: LUT_x0_real_res1 = 121;
            'd122: LUT_x0_real_res1 = 122;
            'd123: LUT_x0_real_res1 = 123;
            'd124: LUT_x0_real_res1 = 124;
            'd125: LUT_x0_real_res1 = 125;
            'd126: LUT_x0_real_res1 = 126;
            'd127: LUT_x0_real_res1 = 127;
            'd128: LUT_x0_real_res1 = 128;
            'd129: LUT_x0_real_res1 = 129;
            'd130: LUT_x0_real_res1 = 130;
            'd131: LUT_x0_real_res1 = 131;
            'd132: LUT_x0_real_res1 = 132;
            'd133: LUT_x0_real_res1 = 133;
            'd134: LUT_x0_real_res1 = 134;
            'd135: LUT_x0_real_res1 = 135;
            'd136: LUT_x0_real_res1 = 136;
            'd137: LUT_x0_real_res1 = 137;
            'd138: LUT_x0_real_res1 = 138;
            'd139: LUT_x0_real_res1 = 139;
            'd140: LUT_x0_real_res1 = 140;
            'd141: LUT_x0_real_res1 = 141;
            'd142: LUT_x0_real_res1 = 142;
            'd143: LUT_x0_real_res1 = 143;
            'd144: LUT_x0_real_res1 = 144;
            'd145: LUT_x0_real_res1 = 145;
            'd146: LUT_x0_real_res1 = 146;
            'd147: LUT_x0_real_res1 = 147;
            'd148: LUT_x0_real_res1 = 148;
            'd149: LUT_x0_real_res1 = 149;
            'd150: LUT_x0_real_res1 = 150;
            'd151: LUT_x0_real_res1 = 151;
            'd152: LUT_x0_real_res1 = 152;
            'd153: LUT_x0_real_res1 = 153;
            'd154: LUT_x0_real_res1 = 154;
            'd155: LUT_x0_real_res1 = 155;
            'd156: LUT_x0_real_res1 = 156;
            'd157: LUT_x0_real_res1 = 157;
            'd158: LUT_x0_real_res1 = 158;
            'd159: LUT_x0_real_res1 = 159;
            'd160: LUT_x0_real_res1 = 160;
            'd161: LUT_x0_real_res1 = 161;
            'd162: LUT_x0_real_res1 = 162;
            'd163: LUT_x0_real_res1 = 163;
            'd164: LUT_x0_real_res1 = 164;
            'd165: LUT_x0_real_res1 = 165;
            'd166: LUT_x0_real_res1 = 166;
            'd167: LUT_x0_real_res1 = 167;
            'd168: LUT_x0_real_res1 = 168;
            'd169: LUT_x0_real_res1 = 169;
            'd170: LUT_x0_real_res1 = 170;
            'd171: LUT_x0_real_res1 = 171;
            'd172: LUT_x0_real_res1 = 172;
            'd173: LUT_x0_real_res1 = 173;
            'd174: LUT_x0_real_res1 = 174;
            'd175: LUT_x0_real_res1 = 175;
            'd176: LUT_x0_real_res1 = 176;
            'd177: LUT_x0_real_res1 = 177;
            'd178: LUT_x0_real_res1 = 178;
            'd179: LUT_x0_real_res1 = 179;
            'd180: LUT_x0_real_res1 = 180;
            'd181: LUT_x0_real_res1 = 181;
            'd182: LUT_x0_real_res1 = 182;
            'd183: LUT_x0_real_res1 = 183;
            'd184: LUT_x0_real_res1 = 184;
            'd185: LUT_x0_real_res1 = 185;
            'd186: LUT_x0_real_res1 = 186;
            'd187: LUT_x0_real_res1 = 187;
            'd188: LUT_x0_real_res1 = 188;
            'd189: LUT_x0_real_res1 = 189;
            'd190: LUT_x0_real_res1 = 190;
            'd191: LUT_x0_real_res1 = 191;
            'd192: LUT_x0_real_res1 = 192;
            'd193: LUT_x0_real_res1 = 193;
            'd194: LUT_x0_real_res1 = 194;
            'd195: LUT_x0_real_res1 = 195;
            'd196: LUT_x0_real_res1 = 196;
            'd197: LUT_x0_real_res1 = 197;
            'd198: LUT_x0_real_res1 = 198;
            'd199: LUT_x0_real_res1 = 199;
            'd200: LUT_x0_real_res1 = 200;
            'd201: LUT_x0_real_res1 = 201;
            'd202: LUT_x0_real_res1 = 202;
            'd203: LUT_x0_real_res1 = 203;
            'd204: LUT_x0_real_res1 = 204;
            'd205: LUT_x0_real_res1 = 205;
            'd206: LUT_x0_real_res1 = 206;
            'd207: LUT_x0_real_res1 = 207;
            'd208: LUT_x0_real_res1 = 208;
            'd209: LUT_x0_real_res1 = 209;
            'd210: LUT_x0_real_res1 = 210;
            'd211: LUT_x0_real_res1 = 211;
            'd212: LUT_x0_real_res1 = 212;
            'd213: LUT_x0_real_res1 = 213;
            'd214: LUT_x0_real_res1 = 214;
            'd215: LUT_x0_real_res1 = 215;
            'd216: LUT_x0_real_res1 = 216;
            'd217: LUT_x0_real_res1 = 217;
            'd218: LUT_x0_real_res1 = 218;
            'd219: LUT_x0_real_res1 = 219;
            'd220: LUT_x0_real_res1 = 220;
            'd221: LUT_x0_real_res1 = 221;
            'd222: LUT_x0_real_res1 = 222;
            'd223: LUT_x0_real_res1 = 223;
            'd224: LUT_x0_real_res1 = 224;
            'd225: LUT_x0_real_res1 = 225;
            'd226: LUT_x0_real_res1 = 226;
            'd227: LUT_x0_real_res1 = 227;
            'd228: LUT_x0_real_res1 = 228;
            'd229: LUT_x0_real_res1 = 229;
            'd230: LUT_x0_real_res1 = 230;
            'd231: LUT_x0_real_res1 = 231;
            'd232: LUT_x0_real_res1 = 232;
            'd233: LUT_x0_real_res1 = 233;
            'd234: LUT_x0_real_res1 = 234;
            'd235: LUT_x0_real_res1 = 235;
            'd236: LUT_x0_real_res1 = 236;
            'd237: LUT_x0_real_res1 = 237;
            'd238: LUT_x0_real_res1 = 238;
            'd239: LUT_x0_real_res1 = 239;
            'd240: LUT_x0_real_res1 = 240;
            'd241: LUT_x0_real_res1 = 241;
            'd242: LUT_x0_real_res1 = 242;
            'd243: LUT_x0_real_res1 = 243;
            'd244: LUT_x0_real_res1 = 244;
            'd245: LUT_x0_real_res1 = 245;
            'd246: LUT_x0_real_res1 = 246;
            'd247: LUT_x0_real_res1 = 247;
            'd248: LUT_x0_real_res1 = 248;
            'd249: LUT_x0_real_res1 = 249;
            'd250: LUT_x0_real_res1 = 250;
            'd251: LUT_x0_real_res1 = 251;
            'd252: LUT_x0_real_res1 = 252;
            'd253: LUT_x0_real_res1 = 253;
            'd254: LUT_x0_real_res1 = 254;
            'd255: LUT_x0_real_res1 = 255;
            'd256: LUT_x0_real_res1 = 256;
            default: LUT_x0_real_res1 = 50;
        endcase
    end //end always
    
    //X0, resonator 1, imaginary 
    always @(*) begin
        case(counter) 
            'd1: LUT_x0_im_res1 = 1;
            'd2: LUT_x0_im_res1 = 2;
            'd3: LUT_x0_im_res1 = 3;
            'd4: LUT_x0_im_res1 = 4;
            'd5: LUT_x0_im_res1 = 5;
            'd6: LUT_x0_im_res1 = 6;
            'd7: LUT_x0_im_res1 = 7;
            'd8: LUT_x0_im_res1 = 8;
            'd9: LUT_x0_im_res1 = 9;
            'd10: LUT_x0_im_res1 = 10;
            'd11: LUT_x0_im_res1 = 11;
            'd12: LUT_x0_im_res1 = 12;
            'd13: LUT_x0_im_res1 = 13;
            'd14: LUT_x0_im_res1 = 14;
            'd15: LUT_x0_im_res1 = 15;
            'd16: LUT_x0_im_res1 = 16;
            'd17: LUT_x0_im_res1 = 17;
            'd18: LUT_x0_im_res1 = 18;
            'd19: LUT_x0_im_res1 = 19;
            'd20: LUT_x0_im_res1 = 20;
            'd21: LUT_x0_im_res1 = 21;
            'd22: LUT_x0_im_res1 = 22;
            'd23: LUT_x0_im_res1 = 23;
            'd24: LUT_x0_im_res1 = 24;
            'd25: LUT_x0_im_res1 = 25;
            'd26: LUT_x0_im_res1 = 26;
            'd27: LUT_x0_im_res1 = 27;
            'd28: LUT_x0_im_res1 = 28;
            'd29: LUT_x0_im_res1 = 29;
            'd30: LUT_x0_im_res1 = 30;
            'd31: LUT_x0_im_res1 = 31;
            'd32: LUT_x0_im_res1 = 32;
            'd33: LUT_x0_im_res1 = 33;
            'd34: LUT_x0_im_res1 = 34;
            'd35: LUT_x0_im_res1 = 35;
            'd36: LUT_x0_im_res1 = 36;
            'd37: LUT_x0_im_res1 = 37;
            'd38: LUT_x0_im_res1 = 38;
            'd39: LUT_x0_im_res1 = 39;
            'd40: LUT_x0_im_res1 = 40;
            'd41: LUT_x0_im_res1 = 41;
            'd42: LUT_x0_im_res1 = 42;
            'd43: LUT_x0_im_res1 = 43;
            'd44: LUT_x0_im_res1 = 44;
            'd45: LUT_x0_im_res1 = 45;
            'd46: LUT_x0_im_res1 = 46;
            'd47: LUT_x0_im_res1 = 47;
            'd48: LUT_x0_im_res1 = 48;
            'd49: LUT_x0_im_res1 = 49;
            'd50: LUT_x0_im_res1 = 50;
            'd51: LUT_x0_im_res1 = 51;
            'd52: LUT_x0_im_res1 = 52;
            'd53: LUT_x0_im_res1 = 53;
            'd54: LUT_x0_im_res1 = 54;
            'd55: LUT_x0_im_res1 = 55;
            'd56: LUT_x0_im_res1 = 56;
            'd57: LUT_x0_im_res1 = 57;
            'd58: LUT_x0_im_res1 = 58;
            'd59: LUT_x0_im_res1 = 59;
            'd60: LUT_x0_im_res1 = 60;
            'd61: LUT_x0_im_res1 = 61;
            'd62: LUT_x0_im_res1 = 62;
            'd63: LUT_x0_im_res1 = 63;
            'd64: LUT_x0_im_res1 = 64;
            'd65: LUT_x0_im_res1 = 65;
            'd66: LUT_x0_im_res1 = 66;
            'd67: LUT_x0_im_res1 = 67;
            'd68: LUT_x0_im_res1 = 68;
            'd69: LUT_x0_im_res1 = 69;
            'd70: LUT_x0_im_res1 = 70;
            'd71: LUT_x0_im_res1 = 71;
            'd72: LUT_x0_im_res1 = 72;
            'd73: LUT_x0_im_res1 = 73;
            'd74: LUT_x0_im_res1 = 74;
            'd75: LUT_x0_im_res1 = 75;
            'd76: LUT_x0_im_res1 = 76;
            'd77: LUT_x0_im_res1 = 77;
            'd78: LUT_x0_im_res1 = 78;
            'd79: LUT_x0_im_res1 = 79;
            'd80: LUT_x0_im_res1 = 80;
            'd81: LUT_x0_im_res1 = 81;
            'd82: LUT_x0_im_res1 = 82;
            'd83: LUT_x0_im_res1 = 83;
            'd84: LUT_x0_im_res1 = 84;
            'd85: LUT_x0_im_res1 = 85;
            'd86: LUT_x0_im_res1 = 86;
            'd87: LUT_x0_im_res1 = 87;
            'd88: LUT_x0_im_res1 = 88;
            'd89: LUT_x0_im_res1 = 89;
            'd90: LUT_x0_im_res1 = 90;
            'd91: LUT_x0_im_res1 = 91;
            'd92: LUT_x0_im_res1 = 92;
            'd93: LUT_x0_im_res1 = 93;
            'd94: LUT_x0_im_res1 = 94;
            'd95: LUT_x0_im_res1 = 95;
            'd96: LUT_x0_im_res1 = 96;
            'd97: LUT_x0_im_res1 = 97;
            'd98: LUT_x0_im_res1 = 98;
            'd99: LUT_x0_im_res1 = 99;
            'd100: LUT_x0_im_res1 = 100;
            'd101: LUT_x0_im_res1 = 101;
            'd102: LUT_x0_im_res1 = 102;
            'd103: LUT_x0_im_res1 = 103;
            'd104: LUT_x0_im_res1 = 104;
            'd105: LUT_x0_im_res1 = 105;
            'd106: LUT_x0_im_res1 = 106;
            'd107: LUT_x0_im_res1 = 107;
            'd108: LUT_x0_im_res1 = 108;
            'd109: LUT_x0_im_res1 = 109;
            'd110: LUT_x0_im_res1 = 110;
            'd111: LUT_x0_im_res1 = 111;
            'd112: LUT_x0_im_res1 = 112;
            'd113: LUT_x0_im_res1 = 113;
            'd114: LUT_x0_im_res1 = 114;
            'd115: LUT_x0_im_res1 = 115;
            'd116: LUT_x0_im_res1 = 116;
            'd117: LUT_x0_im_res1 = 117;
            'd118: LUT_x0_im_res1 = 118;
            'd119: LUT_x0_im_res1 = 119;
            'd120: LUT_x0_im_res1 = 120;
            'd121: LUT_x0_im_res1 = 121;
            'd122: LUT_x0_im_res1 = 122;
            'd123: LUT_x0_im_res1 = 123;
            'd124: LUT_x0_im_res1 = 124;
            'd125: LUT_x0_im_res1 = 125;
            'd126: LUT_x0_im_res1 = 126;
            'd127: LUT_x0_im_res1 = 127;
            'd128: LUT_x0_im_res1 = 128;
            'd129: LUT_x0_im_res1 = 129;
            'd130: LUT_x0_im_res1 = 130;
            'd131: LUT_x0_im_res1 = 131;
            'd132: LUT_x0_im_res1 = 132;
            'd133: LUT_x0_im_res1 = 133;
            'd134: LUT_x0_im_res1 = 134;
            'd135: LUT_x0_im_res1 = 135;
            'd136: LUT_x0_im_res1 = 136;
            'd137: LUT_x0_im_res1 = 137;
            'd138: LUT_x0_im_res1 = 138;
            'd139: LUT_x0_im_res1 = 139;
            'd140: LUT_x0_im_res1 = 140;
            'd141: LUT_x0_im_res1 = 141;
            'd142: LUT_x0_im_res1 = 142;
            'd143: LUT_x0_im_res1 = 143;
            'd144: LUT_x0_im_res1 = 144;
            'd145: LUT_x0_im_res1 = 145;
            'd146: LUT_x0_im_res1 = 146;
            'd147: LUT_x0_im_res1 = 147;
            'd148: LUT_x0_im_res1 = 148;
            'd149: LUT_x0_im_res1 = 149;
            'd150: LUT_x0_im_res1 = 150;
            'd151: LUT_x0_im_res1 = 151;
            'd152: LUT_x0_im_res1 = 152;
            'd153: LUT_x0_im_res1 = 153;
            'd154: LUT_x0_im_res1 = 154;
            'd155: LUT_x0_im_res1 = 155;
            'd156: LUT_x0_im_res1 = 156;
            'd157: LUT_x0_im_res1 = 157;
            'd158: LUT_x0_im_res1 = 158;
            'd159: LUT_x0_im_res1 = 159;
            'd160: LUT_x0_im_res1 = 160;
            'd161: LUT_x0_im_res1 = 161;
            'd162: LUT_x0_im_res1 = 162;
            'd163: LUT_x0_im_res1 = 163;
            'd164: LUT_x0_im_res1 = 164;
            'd165: LUT_x0_im_res1 = 165;
            'd166: LUT_x0_im_res1 = 166;
            'd167: LUT_x0_im_res1 = 167;
            'd168: LUT_x0_im_res1 = 168;
            'd169: LUT_x0_im_res1 = 169;
            'd170: LUT_x0_im_res1 = 170;
            'd171: LUT_x0_im_res1 = 171;
            'd172: LUT_x0_im_res1 = 172;
            'd173: LUT_x0_im_res1 = 173;
            'd174: LUT_x0_im_res1 = 174;
            'd175: LUT_x0_im_res1 = 175;
            'd176: LUT_x0_im_res1 = 176;
            'd177: LUT_x0_im_res1 = 177;
            'd178: LUT_x0_im_res1 = 178;
            'd179: LUT_x0_im_res1 = 179;
            'd180: LUT_x0_im_res1 = 180;
            'd181: LUT_x0_im_res1 = 181;
            'd182: LUT_x0_im_res1 = 182;
            'd183: LUT_x0_im_res1 = 183;
            'd184: LUT_x0_im_res1 = 184;
            'd185: LUT_x0_im_res1 = 185;
            'd186: LUT_x0_im_res1 = 186;
            'd187: LUT_x0_im_res1 = 187;
            'd188: LUT_x0_im_res1 = 188;
            'd189: LUT_x0_im_res1 = 189;
            'd190: LUT_x0_im_res1 = 190;
            'd191: LUT_x0_im_res1 = 191;
            'd192: LUT_x0_im_res1 = 192;
            'd193: LUT_x0_im_res1 = 193;
            'd194: LUT_x0_im_res1 = 194;
            'd195: LUT_x0_im_res1 = 195;
            'd196: LUT_x0_im_res1 = 196;
            'd197: LUT_x0_im_res1 = 197;
            'd198: LUT_x0_im_res1 = 198;
            'd199: LUT_x0_im_res1 = 199;
            'd200: LUT_x0_im_res1 = 200;
            'd201: LUT_x0_im_res1 = 201;
            'd202: LUT_x0_im_res1 = 202;
            'd203: LUT_x0_im_res1 = 203;
            'd204: LUT_x0_im_res1 = 204;
            'd205: LUT_x0_im_res1 = 205;
            'd206: LUT_x0_im_res1 = 206;
            'd207: LUT_x0_im_res1 = 207;
            'd208: LUT_x0_im_res1 = 208;
            'd209: LUT_x0_im_res1 = 209;
            'd210: LUT_x0_im_res1 = 210;
            'd211: LUT_x0_im_res1 = 211;
            'd212: LUT_x0_im_res1 = 212;
            'd213: LUT_x0_im_res1 = 213;
            'd214: LUT_x0_im_res1 = 214;
            'd215: LUT_x0_im_res1 = 215;
            'd216: LUT_x0_im_res1 = 216;
            'd217: LUT_x0_im_res1 = 217;
            'd218: LUT_x0_im_res1 = 218;
            'd219: LUT_x0_im_res1 = 219;
            'd220: LUT_x0_im_res1 = 220;
            'd221: LUT_x0_im_res1 = 221;
            'd222: LUT_x0_im_res1 = 222;
            'd223: LUT_x0_im_res1 = 223;
            'd224: LUT_x0_im_res1 = 224;
            'd225: LUT_x0_im_res1 = 225;
            'd226: LUT_x0_im_res1 = 226;
            'd227: LUT_x0_im_res1 = 227;
            'd228: LUT_x0_im_res1 = 228;
            'd229: LUT_x0_im_res1 = 229;
            'd230: LUT_x0_im_res1 = 230;
            'd231: LUT_x0_im_res1 = 231;
            'd232: LUT_x0_im_res1 = 232;
            'd233: LUT_x0_im_res1 = 233;
            'd234: LUT_x0_im_res1 = 234;
            'd235: LUT_x0_im_res1 = 235;
            'd236: LUT_x0_im_res1 = 236;
            'd237: LUT_x0_im_res1 = 237;
            'd238: LUT_x0_im_res1 = 238;
            'd239: LUT_x0_im_res1 = 239;
            'd240: LUT_x0_im_res1 = 240;
            'd241: LUT_x0_im_res1 = 241;
            'd242: LUT_x0_im_res1 = 242;
            'd243: LUT_x0_im_res1 = 243;
            'd244: LUT_x0_im_res1 = 244;
            'd245: LUT_x0_im_res1 = 245;
            'd246: LUT_x0_im_res1 = 246;
            'd247: LUT_x0_im_res1 = 247;
            'd248: LUT_x0_im_res1 = 248;
            'd249: LUT_x0_im_res1 = 249;
            'd250: LUT_x0_im_res1 = 250;
            'd251: LUT_x0_im_res1 = 251;
            'd252: LUT_x0_im_res1 = 252;
            'd253: LUT_x0_im_res1 = 253;
            'd254: LUT_x0_im_res1 = 254;
            'd255: LUT_x0_im_res1 = 255;
            'd256: LUT_x0_im_res1 = 256;
            default: LUT_x0_im_res1 = 0;
        endcase
    end //end always
    
    //X0, resonator 2, real    
    always @(*) begin
        case(counter) 
            'd1: LUT_x0_real_res2 = 1;
            'd2: LUT_x0_real_res2 = 2;
            'd3: LUT_x0_real_res2 = 3;
            'd4: LUT_x0_real_res2 = 4;
            'd5: LUT_x0_real_res2 = 5;
            'd6: LUT_x0_real_res2 = 6;
            'd7: LUT_x0_real_res2 = 7;
            'd8: LUT_x0_real_res2 = 8;
            'd9: LUT_x0_real_res2 = 9;
            'd10: LUT_x0_real_res2 = 10;
            'd11: LUT_x0_real_res2 = 11;
            'd12: LUT_x0_real_res2 = 12;
            'd13: LUT_x0_real_res2 = 13;
            'd14: LUT_x0_real_res2 = 14;
            'd15: LUT_x0_real_res2 = 15;
            'd16: LUT_x0_real_res2 = 16;
            'd17: LUT_x0_real_res2 = 17;
            'd18: LUT_x0_real_res2 = 18;
            'd19: LUT_x0_real_res2 = 19;
            'd20: LUT_x0_real_res2 = 20;
            'd21: LUT_x0_real_res2 = 21;
            'd22: LUT_x0_real_res2 = 22;
            'd23: LUT_x0_real_res2 = 23;
            'd24: LUT_x0_real_res2 = 24;
            'd25: LUT_x0_real_res2 = 25;
            'd26: LUT_x0_real_res2 = 26;
            'd27: LUT_x0_real_res2 = 27;
            'd28: LUT_x0_real_res2 = 28;
            'd29: LUT_x0_real_res2 = 29;
            'd30: LUT_x0_real_res2 = 30;
            'd31: LUT_x0_real_res2 = 31;
            'd32: LUT_x0_real_res2 = 32;
            'd33: LUT_x0_real_res2 = 33;
            'd34: LUT_x0_real_res2 = 34;
            'd35: LUT_x0_real_res2 = 35;
            'd36: LUT_x0_real_res2 = 36;
            'd37: LUT_x0_real_res2 = 37;
            'd38: LUT_x0_real_res2 = 38;
            'd39: LUT_x0_real_res2 = 39;
            'd40: LUT_x0_real_res2 = 40;
            'd41: LUT_x0_real_res2 = 41;
            'd42: LUT_x0_real_res2 = 42;
            'd43: LUT_x0_real_res2 = 43;
            'd44: LUT_x0_real_res2 = 44;
            'd45: LUT_x0_real_res2 = 45;
            'd46: LUT_x0_real_res2 = 46;
            'd47: LUT_x0_real_res2 = 47;
            'd48: LUT_x0_real_res2 = 48;
            'd49: LUT_x0_real_res2 = 49;
            'd50: LUT_x0_real_res2 = 50;
            'd51: LUT_x0_real_res2 = 51;
            'd52: LUT_x0_real_res2 = 52;
            'd53: LUT_x0_real_res2 = 53;
            'd54: LUT_x0_real_res2 = 54;
            'd55: LUT_x0_real_res2 = 55;
            'd56: LUT_x0_real_res2 = 56;
            'd57: LUT_x0_real_res2 = 57;
            'd58: LUT_x0_real_res2 = 58;
            'd59: LUT_x0_real_res2 = 59;
            'd60: LUT_x0_real_res2 = 60;
            'd61: LUT_x0_real_res2 = 61;
            'd62: LUT_x0_real_res2 = 62;
            'd63: LUT_x0_real_res2 = 63;
            'd64: LUT_x0_real_res2 = 64;
            'd65: LUT_x0_real_res2 = 65;
            'd66: LUT_x0_real_res2 = 66;
            'd67: LUT_x0_real_res2 = 67;
            'd68: LUT_x0_real_res2 = 68;
            'd69: LUT_x0_real_res2 = 69;
            'd70: LUT_x0_real_res2 = 70;
            'd71: LUT_x0_real_res2 = 71;
            'd72: LUT_x0_real_res2 = 72;
            'd73: LUT_x0_real_res2 = 73;
            'd74: LUT_x0_real_res2 = 74;
            'd75: LUT_x0_real_res2 = 75;
            'd76: LUT_x0_real_res2 = 76;
            'd77: LUT_x0_real_res2 = 77;
            'd78: LUT_x0_real_res2 = 78;
            'd79: LUT_x0_real_res2 = 79;
            'd80: LUT_x0_real_res2 = 80;
            'd81: LUT_x0_real_res2 = 81;
            'd82: LUT_x0_real_res2 = 82;
            'd83: LUT_x0_real_res2 = 83;
            'd84: LUT_x0_real_res2 = 84;
            'd85: LUT_x0_real_res2 = 85;
            'd86: LUT_x0_real_res2 = 86;
            'd87: LUT_x0_real_res2 = 87;
            'd88: LUT_x0_real_res2 = 88;
            'd89: LUT_x0_real_res2 = 89;
            'd90: LUT_x0_real_res2 = 90;
            'd91: LUT_x0_real_res2 = 91;
            'd92: LUT_x0_real_res2 = 92;
            'd93: LUT_x0_real_res2 = 93;
            'd94: LUT_x0_real_res2 = 94;
            'd95: LUT_x0_real_res2 = 95;
            'd96: LUT_x0_real_res2 = 96;
            'd97: LUT_x0_real_res2 = 97;
            'd98: LUT_x0_real_res2 = 98;
            'd99: LUT_x0_real_res2 = 99;
            'd100: LUT_x0_real_res2 = 100;
            'd101: LUT_x0_real_res2 = 101;
            'd102: LUT_x0_real_res2 = 102;
            'd103: LUT_x0_real_res2 = 103;
            'd104: LUT_x0_real_res2 = 104;
            'd105: LUT_x0_real_res2 = 105;
            'd106: LUT_x0_real_res2 = 106;
            'd107: LUT_x0_real_res2 = 107;
            'd108: LUT_x0_real_res2 = 108;
            'd109: LUT_x0_real_res2 = 109;
            'd110: LUT_x0_real_res2 = 110;
            'd111: LUT_x0_real_res2 = 111;
            'd112: LUT_x0_real_res2 = 112;
            'd113: LUT_x0_real_res2 = 113;
            'd114: LUT_x0_real_res2 = 114;
            'd115: LUT_x0_real_res2 = 115;
            'd116: LUT_x0_real_res2 = 116;
            'd117: LUT_x0_real_res2 = 117;
            'd118: LUT_x0_real_res2 = 118;
            'd119: LUT_x0_real_res2 = 119;
            'd120: LUT_x0_real_res2 = 120;
            'd121: LUT_x0_real_res2 = 121;
            'd122: LUT_x0_real_res2 = 122;
            'd123: LUT_x0_real_res2 = 123;
            'd124: LUT_x0_real_res2 = 124;
            'd125: LUT_x0_real_res2 = 125;
            'd126: LUT_x0_real_res2 = 126;
            'd127: LUT_x0_real_res2 = 127;
            'd128: LUT_x0_real_res2 = 128;
            'd129: LUT_x0_real_res2 = 129;
            'd130: LUT_x0_real_res2 = 130;
            'd131: LUT_x0_real_res2 = 131;
            'd132: LUT_x0_real_res2 = 132;
            'd133: LUT_x0_real_res2 = 133;
            'd134: LUT_x0_real_res2 = 134;
            'd135: LUT_x0_real_res2 = 135;
            'd136: LUT_x0_real_res2 = 136;
            'd137: LUT_x0_real_res2 = 137;
            'd138: LUT_x0_real_res2 = 138;
            'd139: LUT_x0_real_res2 = 139;
            'd140: LUT_x0_real_res2 = 140;
            'd141: LUT_x0_real_res2 = 141;
            'd142: LUT_x0_real_res2 = 142;
            'd143: LUT_x0_real_res2 = 143;
            'd144: LUT_x0_real_res2 = 144;
            'd145: LUT_x0_real_res2 = 145;
            'd146: LUT_x0_real_res2 = 146;
            'd147: LUT_x0_real_res2 = 147;
            'd148: LUT_x0_real_res2 = 148;
            'd149: LUT_x0_real_res2 = 149;
            'd150: LUT_x0_real_res2 = 150;
            'd151: LUT_x0_real_res2 = 151;
            'd152: LUT_x0_real_res2 = 152;
            'd153: LUT_x0_real_res2 = 153;
            'd154: LUT_x0_real_res2 = 154;
            'd155: LUT_x0_real_res2 = 155;
            'd156: LUT_x0_real_res2 = 156;
            'd157: LUT_x0_real_res2 = 157;
            'd158: LUT_x0_real_res2 = 158;
            'd159: LUT_x0_real_res2 = 159;
            'd160: LUT_x0_real_res2 = 160;
            'd161: LUT_x0_real_res2 = 161;
            'd162: LUT_x0_real_res2 = 162;
            'd163: LUT_x0_real_res2 = 163;
            'd164: LUT_x0_real_res2 = 164;
            'd165: LUT_x0_real_res2 = 165;
            'd166: LUT_x0_real_res2 = 166;
            'd167: LUT_x0_real_res2 = 167;
            'd168: LUT_x0_real_res2 = 168;
            'd169: LUT_x0_real_res2 = 169;
            'd170: LUT_x0_real_res2 = 170;
            'd171: LUT_x0_real_res2 = 171;
            'd172: LUT_x0_real_res2 = 172;
            'd173: LUT_x0_real_res2 = 173;
            'd174: LUT_x0_real_res2 = 174;
            'd175: LUT_x0_real_res2 = 175;
            'd176: LUT_x0_real_res2 = 176;
            'd177: LUT_x0_real_res2 = 177;
            'd178: LUT_x0_real_res2 = 178;
            'd179: LUT_x0_real_res2 = 179;
            'd180: LUT_x0_real_res2 = 180;
            'd181: LUT_x0_real_res2 = 181;
            'd182: LUT_x0_real_res2 = 182;
            'd183: LUT_x0_real_res2 = 183;
            'd184: LUT_x0_real_res2 = 184;
            'd185: LUT_x0_real_res2 = 185;
            'd186: LUT_x0_real_res2 = 186;
            'd187: LUT_x0_real_res2 = 187;
            'd188: LUT_x0_real_res2 = 188;
            'd189: LUT_x0_real_res2 = 189;
            'd190: LUT_x0_real_res2 = 190;
            'd191: LUT_x0_real_res2 = 191;
            'd192: LUT_x0_real_res2 = 192;
            'd193: LUT_x0_real_res2 = 193;
            'd194: LUT_x0_real_res2 = 194;
            'd195: LUT_x0_real_res2 = 195;
            'd196: LUT_x0_real_res2 = 196;
            'd197: LUT_x0_real_res2 = 197;
            'd198: LUT_x0_real_res2 = 198;
            'd199: LUT_x0_real_res2 = 199;
            'd200: LUT_x0_real_res2 = 200;
            'd201: LUT_x0_real_res2 = 201;
            'd202: LUT_x0_real_res2 = 202;
            'd203: LUT_x0_real_res2 = 203;
            'd204: LUT_x0_real_res2 = 204;
            'd205: LUT_x0_real_res2 = 205;
            'd206: LUT_x0_real_res2 = 206;
            'd207: LUT_x0_real_res2 = 207;
            'd208: LUT_x0_real_res2 = 208;
            'd209: LUT_x0_real_res2 = 209;
            'd210: LUT_x0_real_res2 = 210;
            'd211: LUT_x0_real_res2 = 211;
            'd212: LUT_x0_real_res2 = 212;
            'd213: LUT_x0_real_res2 = 213;
            'd214: LUT_x0_real_res2 = 214;
            'd215: LUT_x0_real_res2 = 215;
            'd216: LUT_x0_real_res2 = 216;
            'd217: LUT_x0_real_res2 = 217;
            'd218: LUT_x0_real_res2 = 218;
            'd219: LUT_x0_real_res2 = 219;
            'd220: LUT_x0_real_res2 = 220;
            'd221: LUT_x0_real_res2 = 221;
            'd222: LUT_x0_real_res2 = 222;
            'd223: LUT_x0_real_res2 = 223;
            'd224: LUT_x0_real_res2 = 224;
            'd225: LUT_x0_real_res2 = 225;
            'd226: LUT_x0_real_res2 = 226;
            'd227: LUT_x0_real_res2 = 227;
            'd228: LUT_x0_real_res2 = 228;
            'd229: LUT_x0_real_res2 = 229;
            'd230: LUT_x0_real_res2 = 230;
            'd231: LUT_x0_real_res2 = 231;
            'd232: LUT_x0_real_res2 = 232;
            'd233: LUT_x0_real_res2 = 233;
            'd234: LUT_x0_real_res2 = 234;
            'd235: LUT_x0_real_res2 = 235;
            'd236: LUT_x0_real_res2 = 236;
            'd237: LUT_x0_real_res2 = 237;
            'd238: LUT_x0_real_res2 = 238;
            'd239: LUT_x0_real_res2 = 239;
            'd240: LUT_x0_real_res2 = 240;
            'd241: LUT_x0_real_res2 = 241;
            'd242: LUT_x0_real_res2 = 242;
            'd243: LUT_x0_real_res2 = 243;
            'd244: LUT_x0_real_res2 = 244;
            'd245: LUT_x0_real_res2 = 245;
            'd246: LUT_x0_real_res2 = 246;
            'd247: LUT_x0_real_res2 = 247;
            'd248: LUT_x0_real_res2 = 248;
            'd249: LUT_x0_real_res2 = 249;
            'd250: LUT_x0_real_res2 = 250;
            'd251: LUT_x0_real_res2 = 251;
            'd252: LUT_x0_real_res2 = 252;
            'd253: LUT_x0_real_res2 = 253;
            'd254: LUT_x0_real_res2 = 254;
            'd255: LUT_x0_real_res2 = 255;
            'd256: LUT_x0_real_res2 = 256;
            default: LUT_x0_real_res1 = 0;
        endcase
    end //end always
    
    //X0, resonator 2, imaginary 
    always @(*) begin
        case(counter) 
            'd1: LUT_x0_im_res2 = 1;
            'd2: LUT_x0_im_res2 = 2;
            'd3: LUT_x0_im_res2 = 3;
            'd4: LUT_x0_im_res2 = 4;
            'd5: LUT_x0_im_res2 = 5;
            'd6: LUT_x0_im_res2 = 6;
            'd7: LUT_x0_im_res2 = 7;
            'd8: LUT_x0_im_res2 = 8;
            'd9: LUT_x0_im_res2 = 9;
            'd10: LUT_x0_im_res2 = 10;
            'd11: LUT_x0_im_res2 = 11;
            'd12: LUT_x0_im_res2 = 12;
            'd13: LUT_x0_im_res2 = 13;
            'd14: LUT_x0_im_res2 = 14;
            'd15: LUT_x0_im_res2 = 15;
            'd16: LUT_x0_im_res2 = 16;
            'd17: LUT_x0_im_res2 = 17;
            'd18: LUT_x0_im_res2 = 18;
            'd19: LUT_x0_im_res2 = 19;
            'd20: LUT_x0_im_res2 = 20;
            'd21: LUT_x0_im_res2 = 21;
            'd22: LUT_x0_im_res2 = 22;
            'd23: LUT_x0_im_res2 = 23;
            'd24: LUT_x0_im_res2 = 24;
            'd25: LUT_x0_im_res2 = 25;
            'd26: LUT_x0_im_res2 = 26;
            'd27: LUT_x0_im_res2 = 27;
            'd28: LUT_x0_im_res2 = 28;
            'd29: LUT_x0_im_res2 = 29;
            'd30: LUT_x0_im_res2 = 30;
            'd31: LUT_x0_im_res2 = 31;
            'd32: LUT_x0_im_res2 = 32;
            'd33: LUT_x0_im_res2 = 33;
            'd34: LUT_x0_im_res2 = 34;
            'd35: LUT_x0_im_res2 = 35;
            'd36: LUT_x0_im_res2 = 36;
            'd37: LUT_x0_im_res2 = 37;
            'd38: LUT_x0_im_res2 = 38;
            'd39: LUT_x0_im_res2 = 39;
            'd40: LUT_x0_im_res2 = 40;
            'd41: LUT_x0_im_res2 = 41;
            'd42: LUT_x0_im_res2 = 42;
            'd43: LUT_x0_im_res2 = 43;
            'd44: LUT_x0_im_res2 = 44;
            'd45: LUT_x0_im_res2 = 45;
            'd46: LUT_x0_im_res2 = 46;
            'd47: LUT_x0_im_res2 = 47;
            'd48: LUT_x0_im_res2 = 48;
            'd49: LUT_x0_im_res2 = 49;
            'd50: LUT_x0_im_res2 = 50;
            'd51: LUT_x0_im_res2 = 51;
            'd52: LUT_x0_im_res2 = 52;
            'd53: LUT_x0_im_res2 = 53;
            'd54: LUT_x0_im_res2 = 54;
            'd55: LUT_x0_im_res2 = 55;
            'd56: LUT_x0_im_res2 = 56;
            'd57: LUT_x0_im_res2 = 57;
            'd58: LUT_x0_im_res2 = 58;
            'd59: LUT_x0_im_res2 = 59;
            'd60: LUT_x0_im_res2 = 60;
            'd61: LUT_x0_im_res2 = 61;
            'd62: LUT_x0_im_res2 = 62;
            'd63: LUT_x0_im_res2 = 63;
            'd64: LUT_x0_im_res2 = 64;
            'd65: LUT_x0_im_res2 = 65;
            'd66: LUT_x0_im_res2 = 66;
            'd67: LUT_x0_im_res2 = 67;
            'd68: LUT_x0_im_res2 = 68;
            'd69: LUT_x0_im_res2 = 69;
            'd70: LUT_x0_im_res2 = 70;
            'd71: LUT_x0_im_res2 = 71;
            'd72: LUT_x0_im_res2 = 72;
            'd73: LUT_x0_im_res2 = 73;
            'd74: LUT_x0_im_res2 = 74;
            'd75: LUT_x0_im_res2 = 75;
            'd76: LUT_x0_im_res2 = 76;
            'd77: LUT_x0_im_res2 = 77;
            'd78: LUT_x0_im_res2 = 78;
            'd79: LUT_x0_im_res2 = 79;
            'd80: LUT_x0_im_res2 = 80;
            'd81: LUT_x0_im_res2 = 81;
            'd82: LUT_x0_im_res2 = 82;
            'd83: LUT_x0_im_res2 = 83;
            'd84: LUT_x0_im_res2 = 84;
            'd85: LUT_x0_im_res2 = 85;
            'd86: LUT_x0_im_res2 = 86;
            'd87: LUT_x0_im_res2 = 87;
            'd88: LUT_x0_im_res2 = 88;
            'd89: LUT_x0_im_res2 = 89;
            'd90: LUT_x0_im_res2 = 90;
            'd91: LUT_x0_im_res2 = 91;
            'd92: LUT_x0_im_res2 = 92;
            'd93: LUT_x0_im_res2 = 93;
            'd94: LUT_x0_im_res2 = 94;
            'd95: LUT_x0_im_res2 = 95;
            'd96: LUT_x0_im_res2 = 96;
            'd97: LUT_x0_im_res2 = 97;
            'd98: LUT_x0_im_res2 = 98;
            'd99: LUT_x0_im_res2 = 99;
            'd100: LUT_x0_im_res2 = 100;
            'd101: LUT_x0_im_res2 = 101;
            'd102: LUT_x0_im_res2 = 102;
            'd103: LUT_x0_im_res2 = 103;
            'd104: LUT_x0_im_res2 = 104;
            'd105: LUT_x0_im_res2 = 105;
            'd106: LUT_x0_im_res2 = 106;
            'd107: LUT_x0_im_res2 = 107;
            'd108: LUT_x0_im_res2 = 108;
            'd109: LUT_x0_im_res2 = 109;
            'd110: LUT_x0_im_res2 = 110;
            'd111: LUT_x0_im_res2 = 111;
            'd112: LUT_x0_im_res2 = 112;
            'd113: LUT_x0_im_res2 = 113;
            'd114: LUT_x0_im_res2 = 114;
            'd115: LUT_x0_im_res2 = 115;
            'd116: LUT_x0_im_res2 = 116;
            'd117: LUT_x0_im_res2 = 117;
            'd118: LUT_x0_im_res2 = 118;
            'd119: LUT_x0_im_res2 = 119;
            'd120: LUT_x0_im_res2 = 120;
            'd121: LUT_x0_im_res2 = 121;
            'd122: LUT_x0_im_res2 = 122;
            'd123: LUT_x0_im_res2 = 123;
            'd124: LUT_x0_im_res2 = 124;
            'd125: LUT_x0_im_res2 = 125;
            'd126: LUT_x0_im_res2 = 126;
            'd127: LUT_x0_im_res2 = 127;
            'd128: LUT_x0_im_res2 = 128;
            'd129: LUT_x0_im_res2 = 129;
            'd130: LUT_x0_im_res2 = 130;
            'd131: LUT_x0_im_res2 = 131;
            'd132: LUT_x0_im_res2 = 132;
            'd133: LUT_x0_im_res2 = 133;
            'd134: LUT_x0_im_res2 = 134;
            'd135: LUT_x0_im_res2 = 135;
            'd136: LUT_x0_im_res2 = 136;
            'd137: LUT_x0_im_res2 = 137;
            'd138: LUT_x0_im_res2 = 138;
            'd139: LUT_x0_im_res2 = 139;
            'd140: LUT_x0_im_res2 = 140;
            'd141: LUT_x0_im_res2 = 141;
            'd142: LUT_x0_im_res2 = 142;
            'd143: LUT_x0_im_res2 = 143;
            'd144: LUT_x0_im_res2 = 144;
            'd145: LUT_x0_im_res2 = 145;
            'd146: LUT_x0_im_res2 = 146;
            'd147: LUT_x0_im_res2 = 147;
            'd148: LUT_x0_im_res2 = 148;
            'd149: LUT_x0_im_res2 = 149;
            'd150: LUT_x0_im_res2 = 150;
            'd151: LUT_x0_im_res2 = 151;
            'd152: LUT_x0_im_res2 = 152;
            'd153: LUT_x0_im_res2 = 153;
            'd154: LUT_x0_im_res2 = 154;
            'd155: LUT_x0_im_res2 = 155;
            'd156: LUT_x0_im_res2 = 156;
            'd157: LUT_x0_im_res2 = 157;
            'd158: LUT_x0_im_res2 = 158;
            'd159: LUT_x0_im_res2 = 159;
            'd160: LUT_x0_im_res2 = 160;
            'd161: LUT_x0_im_res2 = 161;
            'd162: LUT_x0_im_res2 = 162;
            'd163: LUT_x0_im_res2 = 163;
            'd164: LUT_x0_im_res2 = 164;
            'd165: LUT_x0_im_res2 = 165;
            'd166: LUT_x0_im_res2 = 166;
            'd167: LUT_x0_im_res2 = 167;
            'd168: LUT_x0_im_res2 = 168;
            'd169: LUT_x0_im_res2 = 169;
            'd170: LUT_x0_im_res2 = 170;
            'd171: LUT_x0_im_res2 = 171;
            'd172: LUT_x0_im_res2 = 172;
            'd173: LUT_x0_im_res2 = 173;
            'd174: LUT_x0_im_res2 = 174;
            'd175: LUT_x0_im_res2 = 175;
            'd176: LUT_x0_im_res2 = 176;
            'd177: LUT_x0_im_res2 = 177;
            'd178: LUT_x0_im_res2 = 178;
            'd179: LUT_x0_im_res2 = 179;
            'd180: LUT_x0_im_res2 = 180;
            'd181: LUT_x0_im_res2 = 181;
            'd182: LUT_x0_im_res2 = 182;
            'd183: LUT_x0_im_res2 = 183;
            'd184: LUT_x0_im_res2 = 184;
            'd185: LUT_x0_im_res2 = 185;
            'd186: LUT_x0_im_res2 = 186;
            'd187: LUT_x0_im_res2 = 187;
            'd188: LUT_x0_im_res2 = 188;
            'd189: LUT_x0_im_res2 = 189;
            'd190: LUT_x0_im_res2 = 190;
            'd191: LUT_x0_im_res2 = 191;
            'd192: LUT_x0_im_res2 = 192;
            'd193: LUT_x0_im_res2 = 193;
            'd194: LUT_x0_im_res2 = 194;
            'd195: LUT_x0_im_res2 = 195;
            'd196: LUT_x0_im_res2 = 196;
            'd197: LUT_x0_im_res2 = 197;
            'd198: LUT_x0_im_res2 = 198;
            'd199: LUT_x0_im_res2 = 199;
            'd200: LUT_x0_im_res2 = 200;
            'd201: LUT_x0_im_res2 = 201;
            'd202: LUT_x0_im_res2 = 202;
            'd203: LUT_x0_im_res2 = 203;
            'd204: LUT_x0_im_res2 = 204;
            'd205: LUT_x0_im_res2 = 205;
            'd206: LUT_x0_im_res2 = 206;
            'd207: LUT_x0_im_res2 = 207;
            'd208: LUT_x0_im_res2 = 208;
            'd209: LUT_x0_im_res2 = 209;
            'd210: LUT_x0_im_res2 = 210;
            'd211: LUT_x0_im_res2 = 211;
            'd212: LUT_x0_im_res2 = 212;
            'd213: LUT_x0_im_res2 = 213;
            'd214: LUT_x0_im_res2 = 214;
            'd215: LUT_x0_im_res2 = 215;
            'd216: LUT_x0_im_res2 = 216;
            'd217: LUT_x0_im_res2 = 217;
            'd218: LUT_x0_im_res2 = 218;
            'd219: LUT_x0_im_res2 = 219;
            'd220: LUT_x0_im_res2 = 220;
            'd221: LUT_x0_im_res2 = 221;
            'd222: LUT_x0_im_res2 = 222;
            'd223: LUT_x0_im_res2 = 223;
            'd224: LUT_x0_im_res2 = 224;
            'd225: LUT_x0_im_res2 = 225;
            'd226: LUT_x0_im_res2 = 226;
            'd227: LUT_x0_im_res2 = 227;
            'd228: LUT_x0_im_res2 = 228;
            'd229: LUT_x0_im_res2 = 229;
            'd230: LUT_x0_im_res2 = 230;
            'd231: LUT_x0_im_res2 = 231;
            'd232: LUT_x0_im_res2 = 232;
            'd233: LUT_x0_im_res2 = 233;
            'd234: LUT_x0_im_res2 = 234;
            'd235: LUT_x0_im_res2 = 235;
            'd236: LUT_x0_im_res2 = 236;
            'd237: LUT_x0_im_res2 = 237;
            'd238: LUT_x0_im_res2 = 238;
            'd239: LUT_x0_im_res2 = 239;
            'd240: LUT_x0_im_res2 = 240;
            'd241: LUT_x0_im_res2 = 241;
            'd242: LUT_x0_im_res2 = 242;
            'd243: LUT_x0_im_res2 = 243;
            'd244: LUT_x0_im_res2 = 244;
            'd245: LUT_x0_im_res2 = 245;
            'd246: LUT_x0_im_res2 = 246;
            'd247: LUT_x0_im_res2 = 247;
            'd248: LUT_x0_im_res2 = 248;
            'd249: LUT_x0_im_res2 = 249;
            'd250: LUT_x0_im_res2 = 250;
            'd251: LUT_x0_im_res2 = 251;
            'd252: LUT_x0_im_res2 = 252;
            'd253: LUT_x0_im_res2 = 253;
            'd254: LUT_x0_im_res2 = 254;
            'd255: LUT_x0_im_res2 = 255;
            'd256: LUT_x0_im_res2 = 256;
            default: LUT_x0_im_res1 = 0;
        endcase
    end //end always

    
    //X1, resonator 1, real    
    always @(*) begin
        case(counter) 
            'd1: LUT_x1_real_res1 = 1;
            'd2: LUT_x1_real_res1 = 2;
            'd3: LUT_x1_real_res1 = 3;
            'd4: LUT_x1_real_res1 = 4;
            'd5: LUT_x1_real_res1 = 5;
            'd6: LUT_x1_real_res1 = 6;
            'd7: LUT_x1_real_res1 = 7;
            'd8: LUT_x1_real_res1 = 8;
            'd9: LUT_x1_real_res1 = 9;
            'd10: LUT_x1_real_res1 = 10;
            'd11: LUT_x1_real_res1 = 11;
            'd12: LUT_x1_real_res1 = 12;
            'd13: LUT_x1_real_res1 = 13;
            'd14: LUT_x1_real_res1 = 14;
            'd15: LUT_x1_real_res1 = 15;
            'd16: LUT_x1_real_res1 = 16;
            'd17: LUT_x1_real_res1 = 17;
            'd18: LUT_x1_real_res1 = 18;
            'd19: LUT_x1_real_res1 = 19;
            'd20: LUT_x1_real_res1 = 20;
            'd21: LUT_x1_real_res1 = 21;
            'd22: LUT_x1_real_res1 = 22;
            'd23: LUT_x1_real_res1 = 23;
            'd24: LUT_x1_real_res1 = 24;
            'd25: LUT_x1_real_res1 = 25;
            'd26: LUT_x1_real_res1 = 26;
            'd27: LUT_x1_real_res1 = 27;
            'd28: LUT_x1_real_res1 = 28;
            'd29: LUT_x1_real_res1 = 29;
            'd30: LUT_x1_real_res1 = 30;
            'd31: LUT_x1_real_res1 = 31;
            'd32: LUT_x1_real_res1 = 32;
            'd33: LUT_x1_real_res1 = 33;
            'd34: LUT_x1_real_res1 = 34;
            'd35: LUT_x1_real_res1 = 35;
            'd36: LUT_x1_real_res1 = 36;
            'd37: LUT_x1_real_res1 = 37;
            'd38: LUT_x1_real_res1 = 38;
            'd39: LUT_x1_real_res1 = 39;
            'd40: LUT_x1_real_res1 = 40;
            'd41: LUT_x1_real_res1 = 41;
            'd42: LUT_x1_real_res1 = 42;
            'd43: LUT_x1_real_res1 = 43;
            'd44: LUT_x1_real_res1 = 44;
            'd45: LUT_x1_real_res1 = 45;
            'd46: LUT_x1_real_res1 = 46;
            'd47: LUT_x1_real_res1 = 47;
            'd48: LUT_x1_real_res1 = 48;
            'd49: LUT_x1_real_res1 = 49;
            'd50: LUT_x1_real_res1 = 50;
            'd51: LUT_x1_real_res1 = 51;
            'd52: LUT_x1_real_res1 = 52;
            'd53: LUT_x1_real_res1 = 53;
            'd54: LUT_x1_real_res1 = 54;
            'd55: LUT_x1_real_res1 = 55;
            'd56: LUT_x1_real_res1 = 56;
            'd57: LUT_x1_real_res1 = 57;
            'd58: LUT_x1_real_res1 = 58;
            'd59: LUT_x1_real_res1 = 59;
            'd60: LUT_x1_real_res1 = 60;
            'd61: LUT_x1_real_res1 = 61;
            'd62: LUT_x1_real_res1 = 62;
            'd63: LUT_x1_real_res1 = 63;
            'd64: LUT_x1_real_res1 = 64;
            'd65: LUT_x1_real_res1 = 65;
            'd66: LUT_x1_real_res1 = 66;
            'd67: LUT_x1_real_res1 = 67;
            'd68: LUT_x1_real_res1 = 68;
            'd69: LUT_x1_real_res1 = 69;
            'd70: LUT_x1_real_res1 = 70;
            'd71: LUT_x1_real_res1 = 71;
            'd72: LUT_x1_real_res1 = 72;
            'd73: LUT_x1_real_res1 = 73;
            'd74: LUT_x1_real_res1 = 74;
            'd75: LUT_x1_real_res1 = 75;
            'd76: LUT_x1_real_res1 = 76;
            'd77: LUT_x1_real_res1 = 77;
            'd78: LUT_x1_real_res1 = 78;
            'd79: LUT_x1_real_res1 = 79;
            'd80: LUT_x1_real_res1 = 80;
            'd81: LUT_x1_real_res1 = 81;
            'd82: LUT_x1_real_res1 = 82;
            'd83: LUT_x1_real_res1 = 83;
            'd84: LUT_x1_real_res1 = 84;
            'd85: LUT_x1_real_res1 = 85;
            'd86: LUT_x1_real_res1 = 86;
            'd87: LUT_x1_real_res1 = 87;
            'd88: LUT_x1_real_res1 = 88;
            'd89: LUT_x1_real_res1 = 89;
            'd90: LUT_x1_real_res1 = 90;
            'd91: LUT_x1_real_res1 = 91;
            'd92: LUT_x1_real_res1 = 92;
            'd93: LUT_x1_real_res1 = 93;
            'd94: LUT_x1_real_res1 = 94;
            'd95: LUT_x1_real_res1 = 95;
            'd96: LUT_x1_real_res1 = 96;
            'd97: LUT_x1_real_res1 = 97;
            'd98: LUT_x1_real_res1 = 98;
            'd99: LUT_x1_real_res1 = 99;
            'd100: LUT_x1_real_res1 = 100;
            'd101: LUT_x1_real_res1 = 101;
            'd102: LUT_x1_real_res1 = 102;
            'd103: LUT_x1_real_res1 = 103;
            'd104: LUT_x1_real_res1 = 104;
            'd105: LUT_x1_real_res1 = 105;
            'd106: LUT_x1_real_res1 = 106;
            'd107: LUT_x1_real_res1 = 107;
            'd108: LUT_x1_real_res1 = 108;
            'd109: LUT_x1_real_res1 = 109;
            'd110: LUT_x1_real_res1 = 110;
            'd111: LUT_x1_real_res1 = 111;
            'd112: LUT_x1_real_res1 = 112;
            'd113: LUT_x1_real_res1 = 113;
            'd114: LUT_x1_real_res1 = 114;
            'd115: LUT_x1_real_res1 = 115;
            'd116: LUT_x1_real_res1 = 116;
            'd117: LUT_x1_real_res1 = 117;
            'd118: LUT_x1_real_res1 = 118;
            'd119: LUT_x1_real_res1 = 119;
            'd120: LUT_x1_real_res1 = 120;
            'd121: LUT_x1_real_res1 = 121;
            'd122: LUT_x1_real_res1 = 122;
            'd123: LUT_x1_real_res1 = 123;
            'd124: LUT_x1_real_res1 = 124;
            'd125: LUT_x1_real_res1 = 125;
            'd126: LUT_x1_real_res1 = 126;
            'd127: LUT_x1_real_res1 = 127;
            'd128: LUT_x1_real_res1 = 128;
            'd129: LUT_x1_real_res1 = 129;
            'd130: LUT_x1_real_res1 = 130;
            'd131: LUT_x1_real_res1 = 131;
            'd132: LUT_x1_real_res1 = 132;
            'd133: LUT_x1_real_res1 = 133;
            'd134: LUT_x1_real_res1 = 134;
            'd135: LUT_x1_real_res1 = 135;
            'd136: LUT_x1_real_res1 = 136;
            'd137: LUT_x1_real_res1 = 137;
            'd138: LUT_x1_real_res1 = 138;
            'd139: LUT_x1_real_res1 = 139;
            'd140: LUT_x1_real_res1 = 140;
            'd141: LUT_x1_real_res1 = 141;
            'd142: LUT_x1_real_res1 = 142;
            'd143: LUT_x1_real_res1 = 143;
            'd144: LUT_x1_real_res1 = 144;
            'd145: LUT_x1_real_res1 = 145;
            'd146: LUT_x1_real_res1 = 146;
            'd147: LUT_x1_real_res1 = 147;
            'd148: LUT_x1_real_res1 = 148;
            'd149: LUT_x1_real_res1 = 149;
            'd150: LUT_x1_real_res1 = 150;
            'd151: LUT_x1_real_res1 = 151;
            'd152: LUT_x1_real_res1 = 152;
            'd153: LUT_x1_real_res1 = 153;
            'd154: LUT_x1_real_res1 = 154;
            'd155: LUT_x1_real_res1 = 155;
            'd156: LUT_x1_real_res1 = 156;
            'd157: LUT_x1_real_res1 = 157;
            'd158: LUT_x1_real_res1 = 158;
            'd159: LUT_x1_real_res1 = 159;
            'd160: LUT_x1_real_res1 = 160;
            'd161: LUT_x1_real_res1 = 161;
            'd162: LUT_x1_real_res1 = 162;
            'd163: LUT_x1_real_res1 = 163;
            'd164: LUT_x1_real_res1 = 164;
            'd165: LUT_x1_real_res1 = 165;
            'd166: LUT_x1_real_res1 = 166;
            'd167: LUT_x1_real_res1 = 167;
            'd168: LUT_x1_real_res1 = 168;
            'd169: LUT_x1_real_res1 = 169;
            'd170: LUT_x1_real_res1 = 170;
            'd171: LUT_x1_real_res1 = 171;
            'd172: LUT_x1_real_res1 = 172;
            'd173: LUT_x1_real_res1 = 173;
            'd174: LUT_x1_real_res1 = 174;
            'd175: LUT_x1_real_res1 = 175;
            'd176: LUT_x1_real_res1 = 176;
            'd177: LUT_x1_real_res1 = 177;
            'd178: LUT_x1_real_res1 = 178;
            'd179: LUT_x1_real_res1 = 179;
            'd180: LUT_x1_real_res1 = 180;
            'd181: LUT_x1_real_res1 = 181;
            'd182: LUT_x1_real_res1 = 182;
            'd183: LUT_x1_real_res1 = 183;
            'd184: LUT_x1_real_res1 = 184;
            'd185: LUT_x1_real_res1 = 185;
            'd186: LUT_x1_real_res1 = 186;
            'd187: LUT_x1_real_res1 = 187;
            'd188: LUT_x1_real_res1 = 188;
            'd189: LUT_x1_real_res1 = 189;
            'd190: LUT_x1_real_res1 = 190;
            'd191: LUT_x1_real_res1 = 191;
            'd192: LUT_x1_real_res1 = 192;
            'd193: LUT_x1_real_res1 = 193;
            'd194: LUT_x1_real_res1 = 194;
            'd195: LUT_x1_real_res1 = 195;
            'd196: LUT_x1_real_res1 = 196;
            'd197: LUT_x1_real_res1 = 197;
            'd198: LUT_x1_real_res1 = 198;
            'd199: LUT_x1_real_res1 = 199;
            'd200: LUT_x1_real_res1 = 200;
            'd201: LUT_x1_real_res1 = 201;
            'd202: LUT_x1_real_res1 = 202;
            'd203: LUT_x1_real_res1 = 203;
            'd204: LUT_x1_real_res1 = 204;
            'd205: LUT_x1_real_res1 = 205;
            'd206: LUT_x1_real_res1 = 206;
            'd207: LUT_x1_real_res1 = 207;
            'd208: LUT_x1_real_res1 = 208;
            'd209: LUT_x1_real_res1 = 209;
            'd210: LUT_x1_real_res1 = 210;
            'd211: LUT_x1_real_res1 = 211;
            'd212: LUT_x1_real_res1 = 212;
            'd213: LUT_x1_real_res1 = 213;
            'd214: LUT_x1_real_res1 = 214;
            'd215: LUT_x1_real_res1 = 215;
            'd216: LUT_x1_real_res1 = 216;
            'd217: LUT_x1_real_res1 = 217;
            'd218: LUT_x1_real_res1 = 218;
            'd219: LUT_x1_real_res1 = 219;
            'd220: LUT_x1_real_res1 = 220;
            'd221: LUT_x1_real_res1 = 221;
            'd222: LUT_x1_real_res1 = 222;
            'd223: LUT_x1_real_res1 = 223;
            'd224: LUT_x1_real_res1 = 224;
            'd225: LUT_x1_real_res1 = 225;
            'd226: LUT_x1_real_res1 = 226;
            'd227: LUT_x1_real_res1 = 227;
            'd228: LUT_x1_real_res1 = 228;
            'd229: LUT_x1_real_res1 = 229;
            'd230: LUT_x1_real_res1 = 230;
            'd231: LUT_x1_real_res1 = 231;
            'd232: LUT_x1_real_res1 = 232;
            'd233: LUT_x1_real_res1 = 233;
            'd234: LUT_x1_real_res1 = 234;
            'd235: LUT_x1_real_res1 = 235;
            'd236: LUT_x1_real_res1 = 236;
            'd237: LUT_x1_real_res1 = 237;
            'd238: LUT_x1_real_res1 = 238;
            'd239: LUT_x1_real_res1 = 239;
            'd240: LUT_x1_real_res1 = 240;
            'd241: LUT_x1_real_res1 = 241;
            'd242: LUT_x1_real_res1 = 242;
            'd243: LUT_x1_real_res1 = 243;
            'd244: LUT_x1_real_res1 = 244;
            'd245: LUT_x1_real_res1 = 245;
            'd246: LUT_x1_real_res1 = 246;
            'd247: LUT_x1_real_res1 = 247;
            'd248: LUT_x1_real_res1 = 248;
            'd249: LUT_x1_real_res1 = 249;
            'd250: LUT_x1_real_res1 = 250;
            'd251: LUT_x1_real_res1 = 251;
            'd252: LUT_x1_real_res1 = 252;
            'd253: LUT_x1_real_res1 = 253;
            'd254: LUT_x1_real_res1 = 254;
            'd255: LUT_x1_real_res1 = 255;
            'd256: LUT_x1_real_res1 = 256; 
            default: LUT_x1_real_res1 = 0;
        endcase
    end //end always
    
    //X1, resonator 1, imaginary 
    always @(*) begin
        case(counter) 
            'd1: LUT_x1_im_res1 = 1;
            'd2: LUT_x1_im_res1 = 2;
            'd3: LUT_x1_im_res1 = 3;
            'd4: LUT_x1_im_res1 = 4;
            'd5: LUT_x1_im_res1 = 5;
            'd6: LUT_x1_im_res1 = 6;
            'd7: LUT_x1_im_res1 = 7;
            'd8: LUT_x1_im_res1 = 8;
            'd9: LUT_x1_im_res1 = 9;
            'd10: LUT_x1_im_res1 = 10;
            'd11: LUT_x1_im_res1 = 11;
            'd12: LUT_x1_im_res1 = 12;
            'd13: LUT_x1_im_res1 = 13;
            'd14: LUT_x1_im_res1 = 14;
            'd15: LUT_x1_im_res1 = 15;
            'd16: LUT_x1_im_res1 = 16;
            'd17: LUT_x1_im_res1 = 17;
            'd18: LUT_x1_im_res1 = 18;
            'd19: LUT_x1_im_res1 = 19;
            'd20: LUT_x1_im_res1 = 20;
            'd21: LUT_x1_im_res1 = 21;
            'd22: LUT_x1_im_res1 = 22;
            'd23: LUT_x1_im_res1 = 23;
            'd24: LUT_x1_im_res1 = 24;
            'd25: LUT_x1_im_res1 = 25;
            'd26: LUT_x1_im_res1 = 26;
            'd27: LUT_x1_im_res1 = 27;
            'd28: LUT_x1_im_res1 = 28;
            'd29: LUT_x1_im_res1 = 29;
            'd30: LUT_x1_im_res1 = 30;
            'd31: LUT_x1_im_res1 = 31;
            'd32: LUT_x1_im_res1 = 32;
            'd33: LUT_x1_im_res1 = 33;
            'd34: LUT_x1_im_res1 = 34;
            'd35: LUT_x1_im_res1 = 35;
            'd36: LUT_x1_im_res1 = 36;
            'd37: LUT_x1_im_res1 = 37;
            'd38: LUT_x1_im_res1 = 38;
            'd39: LUT_x1_im_res1 = 39;
            'd40: LUT_x1_im_res1 = 40;
            'd41: LUT_x1_im_res1 = 41;
            'd42: LUT_x1_im_res1 = 42;
            'd43: LUT_x1_im_res1 = 43;
            'd44: LUT_x1_im_res1 = 44;
            'd45: LUT_x1_im_res1 = 45;
            'd46: LUT_x1_im_res1 = 46;
            'd47: LUT_x1_im_res1 = 47;
            'd48: LUT_x1_im_res1 = 48;
            'd49: LUT_x1_im_res1 = 49;
            'd50: LUT_x1_im_res1 = 50;
            'd51: LUT_x1_im_res1 = 51;
            'd52: LUT_x1_im_res1 = 52;
            'd53: LUT_x1_im_res1 = 53;
            'd54: LUT_x1_im_res1 = 54;
            'd55: LUT_x1_im_res1 = 55;
            'd56: LUT_x1_im_res1 = 56;
            'd57: LUT_x1_im_res1 = 57;
            'd58: LUT_x1_im_res1 = 58;
            'd59: LUT_x1_im_res1 = 59;
            'd60: LUT_x1_im_res1 = 60;
            'd61: LUT_x1_im_res1 = 61;
            'd62: LUT_x1_im_res1 = 62;
            'd63: LUT_x1_im_res1 = 63;
            'd64: LUT_x1_im_res1 = 64;
            'd65: LUT_x1_im_res1 = 65;
            'd66: LUT_x1_im_res1 = 66;
            'd67: LUT_x1_im_res1 = 67;
            'd68: LUT_x1_im_res1 = 68;
            'd69: LUT_x1_im_res1 = 69;
            'd70: LUT_x1_im_res1 = 70;
            'd71: LUT_x1_im_res1 = 71;
            'd72: LUT_x1_im_res1 = 72;
            'd73: LUT_x1_im_res1 = 73;
            'd74: LUT_x1_im_res1 = 74;
            'd75: LUT_x1_im_res1 = 75;
            'd76: LUT_x1_im_res1 = 76;
            'd77: LUT_x1_im_res1 = 77;
            'd78: LUT_x1_im_res1 = 78;
            'd79: LUT_x1_im_res1 = 79;
            'd80: LUT_x1_im_res1 = 80;
            'd81: LUT_x1_im_res1 = 81;
            'd82: LUT_x1_im_res1 = 82;
            'd83: LUT_x1_im_res1 = 83;
            'd84: LUT_x1_im_res1 = 84;
            'd85: LUT_x1_im_res1 = 85;
            'd86: LUT_x1_im_res1 = 86;
            'd87: LUT_x1_im_res1 = 87;
            'd88: LUT_x1_im_res1 = 88;
            'd89: LUT_x1_im_res1 = 89;
            'd90: LUT_x1_im_res1 = 90;
            'd91: LUT_x1_im_res1 = 91;
            'd92: LUT_x1_im_res1 = 92;
            'd93: LUT_x1_im_res1 = 93;
            'd94: LUT_x1_im_res1 = 94;
            'd95: LUT_x1_im_res1 = 95;
            'd96: LUT_x1_im_res1 = 96;
            'd97: LUT_x1_im_res1 = 97;
            'd98: LUT_x1_im_res1 = 98;
            'd99: LUT_x1_im_res1 = 99;
            'd100: LUT_x1_im_res1 = 100;
            'd101: LUT_x1_im_res1 = 101;
            'd102: LUT_x1_im_res1 = 102;
            'd103: LUT_x1_im_res1 = 103;
            'd104: LUT_x1_im_res1 = 104;
            'd105: LUT_x1_im_res1 = 105;
            'd106: LUT_x1_im_res1 = 106;
            'd107: LUT_x1_im_res1 = 107;
            'd108: LUT_x1_im_res1 = 108;
            'd109: LUT_x1_im_res1 = 109;
            'd110: LUT_x1_im_res1 = 110;
            'd111: LUT_x1_im_res1 = 111;
            'd112: LUT_x1_im_res1 = 112;
            'd113: LUT_x1_im_res1 = 113;
            'd114: LUT_x1_im_res1 = 114;
            'd115: LUT_x1_im_res1 = 115;
            'd116: LUT_x1_im_res1 = 116;
            'd117: LUT_x1_im_res1 = 117;
            'd118: LUT_x1_im_res1 = 118;
            'd119: LUT_x1_im_res1 = 119;
            'd120: LUT_x1_im_res1 = 120;
            'd121: LUT_x1_im_res1 = 121;
            'd122: LUT_x1_im_res1 = 122;
            'd123: LUT_x1_im_res1 = 123;
            'd124: LUT_x1_im_res1 = 124;
            'd125: LUT_x1_im_res1 = 125;
            'd126: LUT_x1_im_res1 = 126;
            'd127: LUT_x1_im_res1 = 127;
            'd128: LUT_x1_im_res1 = 128;
            'd129: LUT_x1_im_res1 = 129;
            'd130: LUT_x1_im_res1 = 130;
            'd131: LUT_x1_im_res1 = 131;
            'd132: LUT_x1_im_res1 = 132;
            'd133: LUT_x1_im_res1 = 133;
            'd134: LUT_x1_im_res1 = 134;
            'd135: LUT_x1_im_res1 = 135;
            'd136: LUT_x1_im_res1 = 136;
            'd137: LUT_x1_im_res1 = 137;
            'd138: LUT_x1_im_res1 = 138;
            'd139: LUT_x1_im_res1 = 139;
            'd140: LUT_x1_im_res1 = 140;
            'd141: LUT_x1_im_res1 = 141;
            'd142: LUT_x1_im_res1 = 142;
            'd143: LUT_x1_im_res1 = 143;
            'd144: LUT_x1_im_res1 = 144;
            'd145: LUT_x1_im_res1 = 145;
            'd146: LUT_x1_im_res1 = 146;
            'd147: LUT_x1_im_res1 = 147;
            'd148: LUT_x1_im_res1 = 148;
            'd149: LUT_x1_im_res1 = 149;
            'd150: LUT_x1_im_res1 = 150;
            'd151: LUT_x1_im_res1 = 151;
            'd152: LUT_x1_im_res1 = 152;
            'd153: LUT_x1_im_res1 = 153;
            'd154: LUT_x1_im_res1 = 154;
            'd155: LUT_x1_im_res1 = 155;
            'd156: LUT_x1_im_res1 = 156;
            'd157: LUT_x1_im_res1 = 157;
            'd158: LUT_x1_im_res1 = 158;
            'd159: LUT_x1_im_res1 = 159;
            'd160: LUT_x1_im_res1 = 160;
            'd161: LUT_x1_im_res1 = 161;
            'd162: LUT_x1_im_res1 = 162;
            'd163: LUT_x1_im_res1 = 163;
            'd164: LUT_x1_im_res1 = 164;
            'd165: LUT_x1_im_res1 = 165;
            'd166: LUT_x1_im_res1 = 166;
            'd167: LUT_x1_im_res1 = 167;
            'd168: LUT_x1_im_res1 = 168;
            'd169: LUT_x1_im_res1 = 169;
            'd170: LUT_x1_im_res1 = 170;
            'd171: LUT_x1_im_res1 = 171;
            'd172: LUT_x1_im_res1 = 172;
            'd173: LUT_x1_im_res1 = 173;
            'd174: LUT_x1_im_res1 = 174;
            'd175: LUT_x1_im_res1 = 175;
            'd176: LUT_x1_im_res1 = 176;
            'd177: LUT_x1_im_res1 = 177;
            'd178: LUT_x1_im_res1 = 178;
            'd179: LUT_x1_im_res1 = 179;
            'd180: LUT_x1_im_res1 = 180;
            'd181: LUT_x1_im_res1 = 181;
            'd182: LUT_x1_im_res1 = 182;
            'd183: LUT_x1_im_res1 = 183;
            'd184: LUT_x1_im_res1 = 184;
            'd185: LUT_x1_im_res1 = 185;
            'd186: LUT_x1_im_res1 = 186;
            'd187: LUT_x1_im_res1 = 187;
            'd188: LUT_x1_im_res1 = 188;
            'd189: LUT_x1_im_res1 = 189;
            'd190: LUT_x1_im_res1 = 190;
            'd191: LUT_x1_im_res1 = 191;
            'd192: LUT_x1_im_res1 = 192;
            'd193: LUT_x1_im_res1 = 193;
            'd194: LUT_x1_im_res1 = 194;
            'd195: LUT_x1_im_res1 = 195;
            'd196: LUT_x1_im_res1 = 196;
            'd197: LUT_x1_im_res1 = 197;
            'd198: LUT_x1_im_res1 = 198;
            'd199: LUT_x1_im_res1 = 199;
            'd200: LUT_x1_im_res1 = 200;
            'd201: LUT_x1_im_res1 = 201;
            'd202: LUT_x1_im_res1 = 202;
            'd203: LUT_x1_im_res1 = 203;
            'd204: LUT_x1_im_res1 = 204;
            'd205: LUT_x1_im_res1 = 205;
            'd206: LUT_x1_im_res1 = 206;
            'd207: LUT_x1_im_res1 = 207;
            'd208: LUT_x1_im_res1 = 208;
            'd209: LUT_x1_im_res1 = 209;
            'd210: LUT_x1_im_res1 = 210;
            'd211: LUT_x1_im_res1 = 211;
            'd212: LUT_x1_im_res1 = 212;
            'd213: LUT_x1_im_res1 = 213;
            'd214: LUT_x1_im_res1 = 214;
            'd215: LUT_x1_im_res1 = 215;
            'd216: LUT_x1_im_res1 = 216;
            'd217: LUT_x1_im_res1 = 217;
            'd218: LUT_x1_im_res1 = 218;
            'd219: LUT_x1_im_res1 = 219;
            'd220: LUT_x1_im_res1 = 220;
            'd221: LUT_x1_im_res1 = 221;
            'd222: LUT_x1_im_res1 = 222;
            'd223: LUT_x1_im_res1 = 223;
            'd224: LUT_x1_im_res1 = 224;
            'd225: LUT_x1_im_res1 = 225;
            'd226: LUT_x1_im_res1 = 226;
            'd227: LUT_x1_im_res1 = 227;
            'd228: LUT_x1_im_res1 = 228;
            'd229: LUT_x1_im_res1 = 229;
            'd230: LUT_x1_im_res1 = 230;
            'd231: LUT_x1_im_res1 = 231;
            'd232: LUT_x1_im_res1 = 232;
            'd233: LUT_x1_im_res1 = 233;
            'd234: LUT_x1_im_res1 = 234;
            'd235: LUT_x1_im_res1 = 235;
            'd236: LUT_x1_im_res1 = 236;
            'd237: LUT_x1_im_res1 = 237;
            'd238: LUT_x1_im_res1 = 238;
            'd239: LUT_x1_im_res1 = 239;
            'd240: LUT_x1_im_res1 = 240;
            'd241: LUT_x1_im_res1 = 241;
            'd242: LUT_x1_im_res1 = 242;
            'd243: LUT_x1_im_res1 = 243;
            'd244: LUT_x1_im_res1 = 244;
            'd245: LUT_x1_im_res1 = 245;
            'd246: LUT_x1_im_res1 = 246;
            'd247: LUT_x1_im_res1 = 247;
            'd248: LUT_x1_im_res1 = 248;
            'd249: LUT_x1_im_res1 = 249;
            'd250: LUT_x1_im_res1 = 250;
            'd251: LUT_x1_im_res1 = 251;
            'd252: LUT_x1_im_res1 = 252;
            'd253: LUT_x1_im_res1 = 253;
            'd254: LUT_x1_im_res1 = 254;
            'd255: LUT_x1_im_res1 = 255;
            'd256: LUT_x1_im_res1 = 256;
            default: LUT_x1_im_res1 = 0;
        endcase
    end //end always
    
    //X1, resonator 2, real    
    always @(*) begin
        case(counter) 
            'd1: LUT_x1_real_res2 = 1;
            'd2: LUT_x1_real_res2 = 2;
            'd3: LUT_x1_real_res2 = 3;
            'd4: LUT_x1_real_res2 = 4;
            'd5: LUT_x1_real_res2 = 5;
            'd6: LUT_x1_real_res2 = 6;
            'd7: LUT_x1_real_res2 = 7;
            'd8: LUT_x1_real_res2 = 8;
            'd9: LUT_x1_real_res2 = 9;
            'd10: LUT_x1_real_res2 = 10;
            'd11: LUT_x1_real_res2 = 11;
            'd12: LUT_x1_real_res2 = 12;
            'd13: LUT_x1_real_res2 = 13;
            'd14: LUT_x1_real_res2 = 14;
            'd15: LUT_x1_real_res2 = 15;
            'd16: LUT_x1_real_res2 = 16;
            'd17: LUT_x1_real_res2 = 17;
            'd18: LUT_x1_real_res2 = 18;
            'd19: LUT_x1_real_res2 = 19;
            'd20: LUT_x1_real_res2 = 20;
            'd21: LUT_x1_real_res2 = 21;
            'd22: LUT_x1_real_res2 = 22;
            'd23: LUT_x1_real_res2 = 23;
            'd24: LUT_x1_real_res2 = 24;
            'd25: LUT_x1_real_res2 = 25;
            'd26: LUT_x1_real_res2 = 26;
            'd27: LUT_x1_real_res2 = 27;
            'd28: LUT_x1_real_res2 = 28;
            'd29: LUT_x1_real_res2 = 29;
            'd30: LUT_x1_real_res2 = 30;
            'd31: LUT_x1_real_res2 = 31;
            'd32: LUT_x1_real_res2 = 32;
            'd33: LUT_x1_real_res2 = 33;
            'd34: LUT_x1_real_res2 = 34;
            'd35: LUT_x1_real_res2 = 35;
            'd36: LUT_x1_real_res2 = 36;
            'd37: LUT_x1_real_res2 = 37;
            'd38: LUT_x1_real_res2 = 38;
            'd39: LUT_x1_real_res2 = 39;
            'd40: LUT_x1_real_res2 = 40;
            'd41: LUT_x1_real_res2 = 41;
            'd42: LUT_x1_real_res2 = 42;
            'd43: LUT_x1_real_res2 = 43;
            'd44: LUT_x1_real_res2 = 44;
            'd45: LUT_x1_real_res2 = 45;
            'd46: LUT_x1_real_res2 = 46;
            'd47: LUT_x1_real_res2 = 47;
            'd48: LUT_x1_real_res2 = 48;
            'd49: LUT_x1_real_res2 = 49;
            'd50: LUT_x1_real_res2 = 50;
            'd51: LUT_x1_real_res2 = 51;
            'd52: LUT_x1_real_res2 = 52;
            'd53: LUT_x1_real_res2 = 53;
            'd54: LUT_x1_real_res2 = 54;
            'd55: LUT_x1_real_res2 = 55;
            'd56: LUT_x1_real_res2 = 56;
            'd57: LUT_x1_real_res2 = 57;
            'd58: LUT_x1_real_res2 = 58;
            'd59: LUT_x1_real_res2 = 59;
            'd60: LUT_x1_real_res2 = 60;
            'd61: LUT_x1_real_res2 = 61;
            'd62: LUT_x1_real_res2 = 62;
            'd63: LUT_x1_real_res2 = 63;
            'd64: LUT_x1_real_res2 = 64;
            'd65: LUT_x1_real_res2 = 65;
            'd66: LUT_x1_real_res2 = 66;
            'd67: LUT_x1_real_res2 = 67;
            'd68: LUT_x1_real_res2 = 68;
            'd69: LUT_x1_real_res2 = 69;
            'd70: LUT_x1_real_res2 = 70;
            'd71: LUT_x1_real_res2 = 71;
            'd72: LUT_x1_real_res2 = 72;
            'd73: LUT_x1_real_res2 = 73;
            'd74: LUT_x1_real_res2 = 74;
            'd75: LUT_x1_real_res2 = 75;
            'd76: LUT_x1_real_res2 = 76;
            'd77: LUT_x1_real_res2 = 77;
            'd78: LUT_x1_real_res2 = 78;
            'd79: LUT_x1_real_res2 = 79;
            'd80: LUT_x1_real_res2 = 80;
            'd81: LUT_x1_real_res2 = 81;
            'd82: LUT_x1_real_res2 = 82;
            'd83: LUT_x1_real_res2 = 83;
            'd84: LUT_x1_real_res2 = 84;
            'd85: LUT_x1_real_res2 = 85;
            'd86: LUT_x1_real_res2 = 86;
            'd87: LUT_x1_real_res2 = 87;
            'd88: LUT_x1_real_res2 = 88;
            'd89: LUT_x1_real_res2 = 89;
            'd90: LUT_x1_real_res2 = 90;
            'd91: LUT_x1_real_res2 = 91;
            'd92: LUT_x1_real_res2 = 92;
            'd93: LUT_x1_real_res2 = 93;
            'd94: LUT_x1_real_res2 = 94;
            'd95: LUT_x1_real_res2 = 95;
            'd96: LUT_x1_real_res2 = 96;
            'd97: LUT_x1_real_res2 = 97;
            'd98: LUT_x1_real_res2 = 98;
            'd99: LUT_x1_real_res2 = 99;
            'd100: LUT_x1_real_res2 = 100;
            'd101: LUT_x1_real_res2 = 101;
            'd102: LUT_x1_real_res2 = 102;
            'd103: LUT_x1_real_res2 = 103;
            'd104: LUT_x1_real_res2 = 104;
            'd105: LUT_x1_real_res2 = 105;
            'd106: LUT_x1_real_res2 = 106;
            'd107: LUT_x1_real_res2 = 107;
            'd108: LUT_x1_real_res2 = 108;
            'd109: LUT_x1_real_res2 = 109;
            'd110: LUT_x1_real_res2 = 110;
            'd111: LUT_x1_real_res2 = 111;
            'd112: LUT_x1_real_res2 = 112;
            'd113: LUT_x1_real_res2 = 113;
            'd114: LUT_x1_real_res2 = 114;
            'd115: LUT_x1_real_res2 = 115;
            'd116: LUT_x1_real_res2 = 116;
            'd117: LUT_x1_real_res2 = 117;
            'd118: LUT_x1_real_res2 = 118;
            'd119: LUT_x1_real_res2 = 119;
            'd120: LUT_x1_real_res2 = 120;
            'd121: LUT_x1_real_res2 = 121;
            'd122: LUT_x1_real_res2 = 122;
            'd123: LUT_x1_real_res2 = 123;
            'd124: LUT_x1_real_res2 = 124;
            'd125: LUT_x1_real_res2 = 125;
            'd126: LUT_x1_real_res2 = 126;
            'd127: LUT_x1_real_res2 = 127;
            'd128: LUT_x1_real_res2 = 128;
            'd129: LUT_x1_real_res2 = 129;
            'd130: LUT_x1_real_res2 = 130;
            'd131: LUT_x1_real_res2 = 131;
            'd132: LUT_x1_real_res2 = 132;
            'd133: LUT_x1_real_res2 = 133;
            'd134: LUT_x1_real_res2 = 134;
            'd135: LUT_x1_real_res2 = 135;
            'd136: LUT_x1_real_res2 = 136;
            'd137: LUT_x1_real_res2 = 137;
            'd138: LUT_x1_real_res2 = 138;
            'd139: LUT_x1_real_res2 = 139;
            'd140: LUT_x1_real_res2 = 140;
            'd141: LUT_x1_real_res2 = 141;
            'd142: LUT_x1_real_res2 = 142;
            'd143: LUT_x1_real_res2 = 143;
            'd144: LUT_x1_real_res2 = 144;
            'd145: LUT_x1_real_res2 = 145;
            'd146: LUT_x1_real_res2 = 146;
            'd147: LUT_x1_real_res2 = 147;
            'd148: LUT_x1_real_res2 = 148;
            'd149: LUT_x1_real_res2 = 149;
            'd150: LUT_x1_real_res2 = 150;
            'd151: LUT_x1_real_res2 = 151;
            'd152: LUT_x1_real_res2 = 152;
            'd153: LUT_x1_real_res2 = 153;
            'd154: LUT_x1_real_res2 = 154;
            'd155: LUT_x1_real_res2 = 155;
            'd156: LUT_x1_real_res2 = 156;
            'd157: LUT_x1_real_res2 = 157;
            'd158: LUT_x1_real_res2 = 158;
            'd159: LUT_x1_real_res2 = 159;
            'd160: LUT_x1_real_res2 = 160;
            'd161: LUT_x1_real_res2 = 161;
            'd162: LUT_x1_real_res2 = 162;
            'd163: LUT_x1_real_res2 = 163;
            'd164: LUT_x1_real_res2 = 164;
            'd165: LUT_x1_real_res2 = 165;
            'd166: LUT_x1_real_res2 = 166;
            'd167: LUT_x1_real_res2 = 167;
            'd168: LUT_x1_real_res2 = 168;
            'd169: LUT_x1_real_res2 = 169;
            'd170: LUT_x1_real_res2 = 170;
            'd171: LUT_x1_real_res2 = 171;
            'd172: LUT_x1_real_res2 = 172;
            'd173: LUT_x1_real_res2 = 173;
            'd174: LUT_x1_real_res2 = 174;
            'd175: LUT_x1_real_res2 = 175;
            'd176: LUT_x1_real_res2 = 176;
            'd177: LUT_x1_real_res2 = 177;
            'd178: LUT_x1_real_res2 = 178;
            'd179: LUT_x1_real_res2 = 179;
            'd180: LUT_x1_real_res2 = 180;
            'd181: LUT_x1_real_res2 = 181;
            'd182: LUT_x1_real_res2 = 182;
            'd183: LUT_x1_real_res2 = 183;
            'd184: LUT_x1_real_res2 = 184;
            'd185: LUT_x1_real_res2 = 185;
            'd186: LUT_x1_real_res2 = 186;
            'd187: LUT_x1_real_res2 = 187;
            'd188: LUT_x1_real_res2 = 188;
            'd189: LUT_x1_real_res2 = 189;
            'd190: LUT_x1_real_res2 = 190;
            'd191: LUT_x1_real_res2 = 191;
            'd192: LUT_x1_real_res2 = 192;
            'd193: LUT_x1_real_res2 = 193;
            'd194: LUT_x1_real_res2 = 194;
            'd195: LUT_x1_real_res2 = 195;
            'd196: LUT_x1_real_res2 = 196;
            'd197: LUT_x1_real_res2 = 197;
            'd198: LUT_x1_real_res2 = 198;
            'd199: LUT_x1_real_res2 = 199;
            'd200: LUT_x1_real_res2 = 200;
            'd201: LUT_x1_real_res2 = 201;
            'd202: LUT_x1_real_res2 = 202;
            'd203: LUT_x1_real_res2 = 203;
            'd204: LUT_x1_real_res2 = 204;
            'd205: LUT_x1_real_res2 = 205;
            'd206: LUT_x1_real_res2 = 206;
            'd207: LUT_x1_real_res2 = 207;
            'd208: LUT_x1_real_res2 = 208;
            'd209: LUT_x1_real_res2 = 209;
            'd210: LUT_x1_real_res2 = 210;
            'd211: LUT_x1_real_res2 = 211;
            'd212: LUT_x1_real_res2 = 212;
            'd213: LUT_x1_real_res2 = 213;
            'd214: LUT_x1_real_res2 = 214;
            'd215: LUT_x1_real_res2 = 215;
            'd216: LUT_x1_real_res2 = 216;
            'd217: LUT_x1_real_res2 = 217;
            'd218: LUT_x1_real_res2 = 218;
            'd219: LUT_x1_real_res2 = 219;
            'd220: LUT_x1_real_res2 = 220;
            'd221: LUT_x1_real_res2 = 221;
            'd222: LUT_x1_real_res2 = 222;
            'd223: LUT_x1_real_res2 = 223;
            'd224: LUT_x1_real_res2 = 224;
            'd225: LUT_x1_real_res2 = 225;
            'd226: LUT_x1_real_res2 = 226;
            'd227: LUT_x1_real_res2 = 227;
            'd228: LUT_x1_real_res2 = 228;
            'd229: LUT_x1_real_res2 = 229;
            'd230: LUT_x1_real_res2 = 230;
            'd231: LUT_x1_real_res2 = 231;
            'd232: LUT_x1_real_res2 = 232;
            'd233: LUT_x1_real_res2 = 233;
            'd234: LUT_x1_real_res2 = 234;
            'd235: LUT_x1_real_res2 = 235;
            'd236: LUT_x1_real_res2 = 236;
            'd237: LUT_x1_real_res2 = 237;
            'd238: LUT_x1_real_res2 = 238;
            'd239: LUT_x1_real_res2 = 239;
            'd240: LUT_x1_real_res2 = 240;
            'd241: LUT_x1_real_res2 = 241;
            'd242: LUT_x1_real_res2 = 242;
            'd243: LUT_x1_real_res2 = 243;
            'd244: LUT_x1_real_res2 = 244;
            'd245: LUT_x1_real_res2 = 245;
            'd246: LUT_x1_real_res2 = 246;
            'd247: LUT_x1_real_res2 = 247;
            'd248: LUT_x1_real_res2 = 248;
            'd249: LUT_x1_real_res2 = 249;
            'd250: LUT_x1_real_res2 = 250;
            'd251: LUT_x1_real_res2 = 251;
            'd252: LUT_x1_real_res2 = 252;
            'd253: LUT_x1_real_res2 = 253;
            'd254: LUT_x1_real_res2 = 254;
            'd255: LUT_x1_real_res2 = 255;
            'd256: LUT_x1_real_res2 = 256;
            default: LUT_x1_real_res2 = 0;
        endcase
    end //end always
    
    //X1, resonator 2, imaginary 
    always @(*) begin
        case(counter) 
            'd1: LUT_x1_im_res2 = 1;
            'd2: LUT_x1_im_res2 = 2;
            'd3: LUT_x1_im_res2 = 3;
            'd4: LUT_x1_im_res2 = 4;
            'd5: LUT_x1_im_res2 = 5;
            'd6: LUT_x1_im_res2 = 6;
            'd7: LUT_x1_im_res2 = 7;
            'd8: LUT_x1_im_res2 = 8;
            'd9: LUT_x1_im_res2 = 9;
            'd10: LUT_x1_im_res2 = 10;
            'd11: LUT_x1_im_res2 = 11;
            'd12: LUT_x1_im_res2 = 12;
            'd13: LUT_x1_im_res2 = 13;
            'd14: LUT_x1_im_res2 = 14;
            'd15: LUT_x1_im_res2 = 15;
            'd16: LUT_x1_im_res2 = 16;
            'd17: LUT_x1_im_res2 = 17;
            'd18: LUT_x1_im_res2 = 18;
            'd19: LUT_x1_im_res2 = 19;
            'd20: LUT_x1_im_res2 = 20;
            'd21: LUT_x1_im_res2 = 21;
            'd22: LUT_x1_im_res2 = 22;
            'd23: LUT_x1_im_res2 = 23;
            'd24: LUT_x1_im_res2 = 24;
            'd25: LUT_x1_im_res2 = 25;
            'd26: LUT_x1_im_res2 = 26;
            'd27: LUT_x1_im_res2 = 27;
            'd28: LUT_x1_im_res2 = 28;
            'd29: LUT_x1_im_res2 = 29;
            'd30: LUT_x1_im_res2 = 30;
            'd31: LUT_x1_im_res2 = 31;
            'd32: LUT_x1_im_res2 = 32;
            'd33: LUT_x1_im_res2 = 33;
            'd34: LUT_x1_im_res2 = 34;
            'd35: LUT_x1_im_res2 = 35;
            'd36: LUT_x1_im_res2 = 36;
            'd37: LUT_x1_im_res2 = 37;
            'd38: LUT_x1_im_res2 = 38;
            'd39: LUT_x1_im_res2 = 39;
            'd40: LUT_x1_im_res2 = 40;
            'd41: LUT_x1_im_res2 = 41;
            'd42: LUT_x1_im_res2 = 42;
            'd43: LUT_x1_im_res2 = 43;
            'd44: LUT_x1_im_res2 = 44;
            'd45: LUT_x1_im_res2 = 45;
            'd46: LUT_x1_im_res2 = 46;
            'd47: LUT_x1_im_res2 = 47;
            'd48: LUT_x1_im_res2 = 48;
            'd49: LUT_x1_im_res2 = 49;
            'd50: LUT_x1_im_res2 = 50;
            'd51: LUT_x1_im_res2 = 51;
            'd52: LUT_x1_im_res2 = 52;
            'd53: LUT_x1_im_res2 = 53;
            'd54: LUT_x1_im_res2 = 54;
            'd55: LUT_x1_im_res2 = 55;
            'd56: LUT_x1_im_res2 = 56;
            'd57: LUT_x1_im_res2 = 57;
            'd58: LUT_x1_im_res2 = 58;
            'd59: LUT_x1_im_res2 = 59;
            'd60: LUT_x1_im_res2 = 60;
            'd61: LUT_x1_im_res2 = 61;
            'd62: LUT_x1_im_res2 = 62;
            'd63: LUT_x1_im_res2 = 63;
            'd64: LUT_x1_im_res2 = 64;
            'd65: LUT_x1_im_res2 = 65;
            'd66: LUT_x1_im_res2 = 66;
            'd67: LUT_x1_im_res2 = 67;
            'd68: LUT_x1_im_res2 = 68;
            'd69: LUT_x1_im_res2 = 69;
            'd70: LUT_x1_im_res2 = 70;
            'd71: LUT_x1_im_res2 = 71;
            'd72: LUT_x1_im_res2 = 72;
            'd73: LUT_x1_im_res2 = 73;
            'd74: LUT_x1_im_res2 = 74;
            'd75: LUT_x1_im_res2 = 75;
            'd76: LUT_x1_im_res2 = 76;
            'd77: LUT_x1_im_res2 = 77;
            'd78: LUT_x1_im_res2 = 78;
            'd79: LUT_x1_im_res2 = 79;
            'd80: LUT_x1_im_res2 = 80;
            'd81: LUT_x1_im_res2 = 81;
            'd82: LUT_x1_im_res2 = 82;
            'd83: LUT_x1_im_res2 = 83;
            'd84: LUT_x1_im_res2 = 84;
            'd85: LUT_x1_im_res2 = 85;
            'd86: LUT_x1_im_res2 = 86;
            'd87: LUT_x1_im_res2 = 87;
            'd88: LUT_x1_im_res2 = 88;
            'd89: LUT_x1_im_res2 = 89;
            'd90: LUT_x1_im_res2 = 90;
            'd91: LUT_x1_im_res2 = 91;
            'd92: LUT_x1_im_res2 = 92;
            'd93: LUT_x1_im_res2 = 93;
            'd94: LUT_x1_im_res2 = 94;
            'd95: LUT_x1_im_res2 = 95;
            'd96: LUT_x1_im_res2 = 96;
            'd97: LUT_x1_im_res2 = 97;
            'd98: LUT_x1_im_res2 = 98;
            'd99: LUT_x1_im_res2 = 99;
            'd100: LUT_x1_im_res2 = 100;
            'd101: LUT_x1_im_res2 = 101;
            'd102: LUT_x1_im_res2 = 102;
            'd103: LUT_x1_im_res2 = 103;
            'd104: LUT_x1_im_res2 = 104;
            'd105: LUT_x1_im_res2 = 105;
            'd106: LUT_x1_im_res2 = 106;
            'd107: LUT_x1_im_res2 = 107;
            'd108: LUT_x1_im_res2 = 108;
            'd109: LUT_x1_im_res2 = 109;
            'd110: LUT_x1_im_res2 = 110;
            'd111: LUT_x1_im_res2 = 111;
            'd112: LUT_x1_im_res2 = 112;
            'd113: LUT_x1_im_res2 = 113;
            'd114: LUT_x1_im_res2 = 114;
            'd115: LUT_x1_im_res2 = 115;
            'd116: LUT_x1_im_res2 = 116;
            'd117: LUT_x1_im_res2 = 117;
            'd118: LUT_x1_im_res2 = 118;
            'd119: LUT_x1_im_res2 = 119;
            'd120: LUT_x1_im_res2 = 120;
            'd121: LUT_x1_im_res2 = 121;
            'd122: LUT_x1_im_res2 = 122;
            'd123: LUT_x1_im_res2 = 123;
            'd124: LUT_x1_im_res2 = 124;
            'd125: LUT_x1_im_res2 = 125;
            'd126: LUT_x1_im_res2 = 126;
            'd127: LUT_x1_im_res2 = 127;
            'd128: LUT_x1_im_res2 = 128;
            'd129: LUT_x1_im_res2 = 129;
            'd130: LUT_x1_im_res2 = 130;
            'd131: LUT_x1_im_res2 = 131;
            'd132: LUT_x1_im_res2 = 132;
            'd133: LUT_x1_im_res2 = 133;
            'd134: LUT_x1_im_res2 = 134;
            'd135: LUT_x1_im_res2 = 135;
            'd136: LUT_x1_im_res2 = 136;
            'd137: LUT_x1_im_res2 = 137;
            'd138: LUT_x1_im_res2 = 138;
            'd139: LUT_x1_im_res2 = 139;
            'd140: LUT_x1_im_res2 = 140;
            'd141: LUT_x1_im_res2 = 141;
            'd142: LUT_x1_im_res2 = 142;
            'd143: LUT_x1_im_res2 = 143;
            'd144: LUT_x1_im_res2 = 144;
            'd145: LUT_x1_im_res2 = 145;
            'd146: LUT_x1_im_res2 = 146;
            'd147: LUT_x1_im_res2 = 147;
            'd148: LUT_x1_im_res2 = 148;
            'd149: LUT_x1_im_res2 = 149;
            'd150: LUT_x1_im_res2 = 150;
            'd151: LUT_x1_im_res2 = 151;
            'd152: LUT_x1_im_res2 = 152;
            'd153: LUT_x1_im_res2 = 153;
            'd154: LUT_x1_im_res2 = 154;
            'd155: LUT_x1_im_res2 = 155;
            'd156: LUT_x1_im_res2 = 156;
            'd157: LUT_x1_im_res2 = 157;
            'd158: LUT_x1_im_res2 = 158;
            'd159: LUT_x1_im_res2 = 159;
            'd160: LUT_x1_im_res2 = 160;
            'd161: LUT_x1_im_res2 = 161;
            'd162: LUT_x1_im_res2 = 162;
            'd163: LUT_x1_im_res2 = 163;
            'd164: LUT_x1_im_res2 = 164;
            'd165: LUT_x1_im_res2 = 165;
            'd166: LUT_x1_im_res2 = 166;
            'd167: LUT_x1_im_res2 = 167;
            'd168: LUT_x1_im_res2 = 168;
            'd169: LUT_x1_im_res2 = 169;
            'd170: LUT_x1_im_res2 = 170;
            'd171: LUT_x1_im_res2 = 171;
            'd172: LUT_x1_im_res2 = 172;
            'd173: LUT_x1_im_res2 = 173;
            'd174: LUT_x1_im_res2 = 174;
            'd175: LUT_x1_im_res2 = 175;
            'd176: LUT_x1_im_res2 = 176;
            'd177: LUT_x1_im_res2 = 177;
            'd178: LUT_x1_im_res2 = 178;
            'd179: LUT_x1_im_res2 = 179;
            'd180: LUT_x1_im_res2 = 180;
            'd181: LUT_x1_im_res2 = 181;
            'd182: LUT_x1_im_res2 = 182;
            'd183: LUT_x1_im_res2 = 183;
            'd184: LUT_x1_im_res2 = 184;
            'd185: LUT_x1_im_res2 = 185;
            'd186: LUT_x1_im_res2 = 186;
            'd187: LUT_x1_im_res2 = 187;
            'd188: LUT_x1_im_res2 = 188;
            'd189: LUT_x1_im_res2 = 189;
            'd190: LUT_x1_im_res2 = 190;
            'd191: LUT_x1_im_res2 = 191;
            'd192: LUT_x1_im_res2 = 192;
            'd193: LUT_x1_im_res2 = 193;
            'd194: LUT_x1_im_res2 = 194;
            'd195: LUT_x1_im_res2 = 195;
            'd196: LUT_x1_im_res2 = 196;
            'd197: LUT_x1_im_res2 = 197;
            'd198: LUT_x1_im_res2 = 198;
            'd199: LUT_x1_im_res2 = 199;
            'd200: LUT_x1_im_res2 = 200;
            'd201: LUT_x1_im_res2 = 201;
            'd202: LUT_x1_im_res2 = 202;
            'd203: LUT_x1_im_res2 = 203;
            'd204: LUT_x1_im_res2 = 204;
            'd205: LUT_x1_im_res2 = 205;
            'd206: LUT_x1_im_res2 = 206;
            'd207: LUT_x1_im_res2 = 207;
            'd208: LUT_x1_im_res2 = 208;
            'd209: LUT_x1_im_res2 = 209;
            'd210: LUT_x1_im_res2 = 210;
            'd211: LUT_x1_im_res2 = 211;
            'd212: LUT_x1_im_res2 = 212;
            'd213: LUT_x1_im_res2 = 213;
            'd214: LUT_x1_im_res2 = 214;
            'd215: LUT_x1_im_res2 = 215;
            'd216: LUT_x1_im_res2 = 216;
            'd217: LUT_x1_im_res2 = 217;
            'd218: LUT_x1_im_res2 = 218;
            'd219: LUT_x1_im_res2 = 219;
            'd220: LUT_x1_im_res2 = 220;
            'd221: LUT_x1_im_res2 = 221;
            'd222: LUT_x1_im_res2 = 222;
            'd223: LUT_x1_im_res2 = 223;
            'd224: LUT_x1_im_res2 = 224;
            'd225: LUT_x1_im_res2 = 225;
            'd226: LUT_x1_im_res2 = 226;
            'd227: LUT_x1_im_res2 = 227;
            'd228: LUT_x1_im_res2 = 228;
            'd229: LUT_x1_im_res2 = 229;
            'd230: LUT_x1_im_res2 = 230;
            'd231: LUT_x1_im_res2 = 231;
            'd232: LUT_x1_im_res2 = 232;
            'd233: LUT_x1_im_res2 = 233;
            'd234: LUT_x1_im_res2 = 234;
            'd235: LUT_x1_im_res2 = 235;
            'd236: LUT_x1_im_res2 = 236;
            'd237: LUT_x1_im_res2 = 237;
            'd238: LUT_x1_im_res2 = 238;
            'd239: LUT_x1_im_res2 = 239;
            'd240: LUT_x1_im_res2 = 240;
            'd241: LUT_x1_im_res2 = 241;
            'd242: LUT_x1_im_res2 = 242;
            'd243: LUT_x1_im_res2 = 243;
            'd244: LUT_x1_im_res2 = 244;
            'd245: LUT_x1_im_res2 = 245;
            'd246: LUT_x1_im_res2 = 246;
            'd247: LUT_x1_im_res2 = 247;
            'd248: LUT_x1_im_res2 = 248;
            'd249: LUT_x1_im_res2 = 249;
            'd250: LUT_x1_im_res2 = 250;
            'd251: LUT_x1_im_res2 = 251;
            'd252: LUT_x1_im_res2 = 252;
            'd253: LUT_x1_im_res2 = 253;
            'd254: LUT_x1_im_res2 = 254;
            'd255: LUT_x1_im_res2 = 255;
            'd256: LUT_x1_im_res2 = 256;
            default: LUT_x1_im_res2 = 0;
        endcase
    end //end always */
    
    //X2, resonator 1, real
    always @(*) begin
        case(counter) 
            'd1: LUT_x2_real_res1 = 1;
            'd2: LUT_x2_real_res1 = 2;
            'd3: LUT_x2_real_res1 = 3;
            'd4: LUT_x2_real_res1 = 4;
            'd5: LUT_x2_real_res1 = 5;
            'd6: LUT_x2_real_res1 = 6;
            'd7: LUT_x2_real_res1 = 7;
            'd8: LUT_x2_real_res1 = 8;
            'd9: LUT_x2_real_res1 = 9;
            'd10: LUT_x2_real_res1 = 10;
            'd11: LUT_x2_real_res1 = 11;
            'd12: LUT_x2_real_res1 = 12;
            'd13: LUT_x2_real_res1 = 13;
            'd14: LUT_x2_real_res1 = 14;
            'd15: LUT_x2_real_res1 = 15;
            'd16: LUT_x2_real_res1 = 16;
            'd17: LUT_x2_real_res1 = 17;
            'd18: LUT_x2_real_res1 = 18;
            'd19: LUT_x2_real_res1 = 19;
            'd20: LUT_x2_real_res1 = 20;
            'd21: LUT_x2_real_res1 = 21;
            'd22: LUT_x2_real_res1 = 22;
            'd23: LUT_x2_real_res1 = 23;
            'd24: LUT_x2_real_res1 = 24;
            'd25: LUT_x2_real_res1 = 25;
            'd26: LUT_x2_real_res1 = 26;
            'd27: LUT_x2_real_res1 = 27;
            'd28: LUT_x2_real_res1 = 28;
            'd29: LUT_x2_real_res1 = 29;
            'd30: LUT_x2_real_res1 = 30;
            'd31: LUT_x2_real_res1 = 31;
            'd32: LUT_x2_real_res1 = 32;
            'd33: LUT_x2_real_res1 = 33;
            'd34: LUT_x2_real_res1 = 34;
            'd35: LUT_x2_real_res1 = 35;
            'd36: LUT_x2_real_res1 = 36;
            'd37: LUT_x2_real_res1 = 37;
            'd38: LUT_x2_real_res1 = 38;
            'd39: LUT_x2_real_res1 = 39;
            'd40: LUT_x2_real_res1 = 40;
            'd41: LUT_x2_real_res1 = 41;
            'd42: LUT_x2_real_res1 = 42;
            'd43: LUT_x2_real_res1 = 43;
            'd44: LUT_x2_real_res1 = 44;
            'd45: LUT_x2_real_res1 = 45;
            'd46: LUT_x2_real_res1 = 46;
            'd47: LUT_x2_real_res1 = 47;
            'd48: LUT_x2_real_res1 = 48;
            'd49: LUT_x2_real_res1 = 49;
            'd50: LUT_x2_real_res1 = 50;
            'd51: LUT_x2_real_res1 = 51;
            'd52: LUT_x2_real_res1 = 52;
            'd53: LUT_x2_real_res1 = 53;
            'd54: LUT_x2_real_res1 = 54;
            'd55: LUT_x2_real_res1 = 55;
            'd56: LUT_x2_real_res1 = 56;
            'd57: LUT_x2_real_res1 = 57;
            'd58: LUT_x2_real_res1 = 58;
            'd59: LUT_x2_real_res1 = 59;
            'd60: LUT_x2_real_res1 = 60;
            'd61: LUT_x2_real_res1 = 61;
            'd62: LUT_x2_real_res1 = 62;
            'd63: LUT_x2_real_res1 = 63;
            'd64: LUT_x2_real_res1 = 64;
            'd65: LUT_x2_real_res1 = 65;
            'd66: LUT_x2_real_res1 = 66;
            'd67: LUT_x2_real_res1 = 67;
            'd68: LUT_x2_real_res1 = 68;
            'd69: LUT_x2_real_res1 = 69;
            'd70: LUT_x2_real_res1 = 70;
            'd71: LUT_x2_real_res1 = 71;
            'd72: LUT_x2_real_res1 = 72;
            'd73: LUT_x2_real_res1 = 73;
            'd74: LUT_x2_real_res1 = 74;
            'd75: LUT_x2_real_res1 = 75;
            'd76: LUT_x2_real_res1 = 76;
            'd77: LUT_x2_real_res1 = 77;
            'd78: LUT_x2_real_res1 = 78;
            'd79: LUT_x2_real_res1 = 79;
            'd80: LUT_x2_real_res1 = 80;
            'd81: LUT_x2_real_res1 = 81;
            'd82: LUT_x2_real_res1 = 82;
            'd83: LUT_x2_real_res1 = 83;
            'd84: LUT_x2_real_res1 = 84;
            'd85: LUT_x2_real_res1 = 85;
            'd86: LUT_x2_real_res1 = 86;
            'd87: LUT_x2_real_res1 = 87;
            'd88: LUT_x2_real_res1 = 88;
            'd89: LUT_x2_real_res1 = 89;
            'd90: LUT_x2_real_res1 = 90;
            'd91: LUT_x2_real_res1 = 91;
            'd92: LUT_x2_real_res1 = 92;
            'd93: LUT_x2_real_res1 = 93;
            'd94: LUT_x2_real_res1 = 94;
            'd95: LUT_x2_real_res1 = 95;
            'd96: LUT_x2_real_res1 = 96;
            'd97: LUT_x2_real_res1 = 97;
            'd98: LUT_x2_real_res1 = 98;
            'd99: LUT_x2_real_res1 = 99;
            'd100: LUT_x2_real_res1 = 100;
            'd101: LUT_x2_real_res1 = 101;
            'd102: LUT_x2_real_res1 = 102;
            'd103: LUT_x2_real_res1 = 103;
            'd104: LUT_x2_real_res1 = 104;
            'd105: LUT_x2_real_res1 = 105;
            'd106: LUT_x2_real_res1 = 106;
            'd107: LUT_x2_real_res1 = 107;
            'd108: LUT_x2_real_res1 = 108;
            'd109: LUT_x2_real_res1 = 109;
            'd110: LUT_x2_real_res1 = 110;
            'd111: LUT_x2_real_res1 = 111;
            'd112: LUT_x2_real_res1 = 112;
            'd113: LUT_x2_real_res1 = 113;
            'd114: LUT_x2_real_res1 = 114;
            'd115: LUT_x2_real_res1 = 115;
            'd116: LUT_x2_real_res1 = 116;
            'd117: LUT_x2_real_res1 = 117;
            'd118: LUT_x2_real_res1 = 118;
            'd119: LUT_x2_real_res1 = 119;
            'd120: LUT_x2_real_res1 = 120;
            'd121: LUT_x2_real_res1 = 121;
            'd122: LUT_x2_real_res1 = 122;
            'd123: LUT_x2_real_res1 = 123;
            'd124: LUT_x2_real_res1 = 124;
            'd125: LUT_x2_real_res1 = 125;
            'd126: LUT_x2_real_res1 = 126;
            'd127: LUT_x2_real_res1 = 127;
            'd128: LUT_x2_real_res1 = 128;
            'd129: LUT_x2_real_res1 = 129;
            'd130: LUT_x2_real_res1 = 130;
            'd131: LUT_x2_real_res1 = 131;
            'd132: LUT_x2_real_res1 = 132;
            'd133: LUT_x2_real_res1 = 133;
            'd134: LUT_x2_real_res1 = 134;
            'd135: LUT_x2_real_res1 = 135;
            'd136: LUT_x2_real_res1 = 136;
            'd137: LUT_x2_real_res1 = 137;
            'd138: LUT_x2_real_res1 = 138;
            'd139: LUT_x2_real_res1 = 139;
            'd140: LUT_x2_real_res1 = 140;
            'd141: LUT_x2_real_res1 = 141;
            'd142: LUT_x2_real_res1 = 142;
            'd143: LUT_x2_real_res1 = 143;
            'd144: LUT_x2_real_res1 = 144;
            'd145: LUT_x2_real_res1 = 145;
            'd146: LUT_x2_real_res1 = 146;
            'd147: LUT_x2_real_res1 = 147;
            'd148: LUT_x2_real_res1 = 148;
            'd149: LUT_x2_real_res1 = 149;
            'd150: LUT_x2_real_res1 = 150;
            'd151: LUT_x2_real_res1 = 151;
            'd152: LUT_x2_real_res1 = 152;
            'd153: LUT_x2_real_res1 = 153;
            'd154: LUT_x2_real_res1 = 154;
            'd155: LUT_x2_real_res1 = 155;
            'd156: LUT_x2_real_res1 = 156;
            'd157: LUT_x2_real_res1 = 157;
            'd158: LUT_x2_real_res1 = 158;
            'd159: LUT_x2_real_res1 = 159;
            'd160: LUT_x2_real_res1 = 160;
            'd161: LUT_x2_real_res1 = 161;
            'd162: LUT_x2_real_res1 = 162;
            'd163: LUT_x2_real_res1 = 163;
            'd164: LUT_x2_real_res1 = 164;
            'd165: LUT_x2_real_res1 = 165;
            'd166: LUT_x2_real_res1 = 166;
            'd167: LUT_x2_real_res1 = 167;
            'd168: LUT_x2_real_res1 = 168;
            'd169: LUT_x2_real_res1 = 169;
            'd170: LUT_x2_real_res1 = 170;
            'd171: LUT_x2_real_res1 = 171;
            'd172: LUT_x2_real_res1 = 172;
            'd173: LUT_x2_real_res1 = 173;
            'd174: LUT_x2_real_res1 = 174;
            'd175: LUT_x2_real_res1 = 175;
            'd176: LUT_x2_real_res1 = 176;
            'd177: LUT_x2_real_res1 = 177;
            'd178: LUT_x2_real_res1 = 178;
            'd179: LUT_x2_real_res1 = 179;
            'd180: LUT_x2_real_res1 = 180;
            'd181: LUT_x2_real_res1 = 181;
            'd182: LUT_x2_real_res1 = 182;
            'd183: LUT_x2_real_res1 = 183;
            'd184: LUT_x2_real_res1 = 184;
            'd185: LUT_x2_real_res1 = 185;
            'd186: LUT_x2_real_res1 = 186;
            'd187: LUT_x2_real_res1 = 187;
            'd188: LUT_x2_real_res1 = 188;
            'd189: LUT_x2_real_res1 = 189;
            'd190: LUT_x2_real_res1 = 190;
            'd191: LUT_x2_real_res1 = 191;
            'd192: LUT_x2_real_res1 = 192;
            'd193: LUT_x2_real_res1 = 193;
            'd194: LUT_x2_real_res1 = 194;
            'd195: LUT_x2_real_res1 = 195;
            'd196: LUT_x2_real_res1 = 196;
            'd197: LUT_x2_real_res1 = 197;
            'd198: LUT_x2_real_res1 = 198;
            'd199: LUT_x2_real_res1 = 199;
            'd200: LUT_x2_real_res1 = 200;
            'd201: LUT_x2_real_res1 = 201;
            'd202: LUT_x2_real_res1 = 202;
            'd203: LUT_x2_real_res1 = 203;
            'd204: LUT_x2_real_res1 = 204;
            'd205: LUT_x2_real_res1 = 205;
            'd206: LUT_x2_real_res1 = 206;
            'd207: LUT_x2_real_res1 = 207;
            'd208: LUT_x2_real_res1 = 208;
            'd209: LUT_x2_real_res1 = 209;
            'd210: LUT_x2_real_res1 = 210;
            'd211: LUT_x2_real_res1 = 211;
            'd212: LUT_x2_real_res1 = 212;
            'd213: LUT_x2_real_res1 = 213;
            'd214: LUT_x2_real_res1 = 214;
            'd215: LUT_x2_real_res1 = 215;
            'd216: LUT_x2_real_res1 = 216;
            'd217: LUT_x2_real_res1 = 217;
            'd218: LUT_x2_real_res1 = 218;
            'd219: LUT_x2_real_res1 = 219;
            'd220: LUT_x2_real_res1 = 220;
            'd221: LUT_x2_real_res1 = 221;
            'd222: LUT_x2_real_res1 = 222;
            'd223: LUT_x2_real_res1 = 223;
            'd224: LUT_x2_real_res1 = 224;
            'd225: LUT_x2_real_res1 = 225;
            'd226: LUT_x2_real_res1 = 226;
            'd227: LUT_x2_real_res1 = 227;
            'd228: LUT_x2_real_res1 = 228;
            'd229: LUT_x2_real_res1 = 229;
            'd230: LUT_x2_real_res1 = 230;
            'd231: LUT_x2_real_res1 = 231;
            'd232: LUT_x2_real_res1 = 232;
            'd233: LUT_x2_real_res1 = 233;
            'd234: LUT_x2_real_res1 = 234;
            'd235: LUT_x2_real_res1 = 235;
            'd236: LUT_x2_real_res1 = 236;
            'd237: LUT_x2_real_res1 = 237;
            'd238: LUT_x2_real_res1 = 238;
            'd239: LUT_x2_real_res1 = 239;
            'd240: LUT_x2_real_res1 = 240;
            'd241: LUT_x2_real_res1 = 241;
            'd242: LUT_x2_real_res1 = 242;
            'd243: LUT_x2_real_res1 = 243;
            'd244: LUT_x2_real_res1 = 244;
            'd245: LUT_x2_real_res1 = 245;
            'd246: LUT_x2_real_res1 = 246;
            'd247: LUT_x2_real_res1 = 247;
            'd248: LUT_x2_real_res1 = 248;
            'd249: LUT_x2_real_res1 = 249;
            'd250: LUT_x2_real_res1 = 250;
            'd251: LUT_x2_real_res1 = 251;
            'd252: LUT_x2_real_res1 = 252;
            'd253: LUT_x2_real_res1 = 253;
            'd254: LUT_x2_real_res1 = 254;
            'd255: LUT_x2_real_res1 = 255;
            'd256: LUT_x2_real_res1 = 256;
            default: LUT_x2_real_res1 = 0;
        endcase
    end //end always */
    
    //X2, resonator 1, imaginary
    always @(*) begin
        case(counter) 
            'd1: LUT_x2_im_res1 = 1;
            'd2: LUT_x2_im_res1 = 2;
            'd3: LUT_x2_im_res1 = 3;
            'd4: LUT_x2_im_res1 = 4;
            'd5: LUT_x2_im_res1 = 5;
            'd6: LUT_x2_im_res1 = 6;
            'd7: LUT_x2_im_res1 = 7;
            'd8: LUT_x2_im_res1 = 8;
            'd9: LUT_x2_im_res1 = 9;
            'd10: LUT_x2_im_res1 = 10;
            'd11: LUT_x2_im_res1 = 11;
            'd12: LUT_x2_im_res1 = 12;
            'd13: LUT_x2_im_res1 = 13;
            'd14: LUT_x2_im_res1 = 14;
            'd15: LUT_x2_im_res1 = 15;
            'd16: LUT_x2_im_res1 = 16;
            'd17: LUT_x2_im_res1 = 17;
            'd18: LUT_x2_im_res1 = 18;
            'd19: LUT_x2_im_res1 = 19;
            'd20: LUT_x2_im_res1 = 20;
            'd21: LUT_x2_im_res1 = 21;
            'd22: LUT_x2_im_res1 = 22;
            'd23: LUT_x2_im_res1 = 23;
            'd24: LUT_x2_im_res1 = 24;
            'd25: LUT_x2_im_res1 = 25;
            'd26: LUT_x2_im_res1 = 26;
            'd27: LUT_x2_im_res1 = 27;
            'd28: LUT_x2_im_res1 = 28;
            'd29: LUT_x2_im_res1 = 29;
            'd30: LUT_x2_im_res1 = 30;
            'd31: LUT_x2_im_res1 = 31;
            'd32: LUT_x2_im_res1 = 32;
            'd33: LUT_x2_im_res1 = 33;
            'd34: LUT_x2_im_res1 = 34;
            'd35: LUT_x2_im_res1 = 35;
            'd36: LUT_x2_im_res1 = 36;
            'd37: LUT_x2_im_res1 = 37;
            'd38: LUT_x2_im_res1 = 38;
            'd39: LUT_x2_im_res1 = 39;
            'd40: LUT_x2_im_res1 = 40;
            'd41: LUT_x2_im_res1 = 41;
            'd42: LUT_x2_im_res1 = 42;
            'd43: LUT_x2_im_res1 = 43;
            'd44: LUT_x2_im_res1 = 44;
            'd45: LUT_x2_im_res1 = 45;
            'd46: LUT_x2_im_res1 = 46;
            'd47: LUT_x2_im_res1 = 47;
            'd48: LUT_x2_im_res1 = 48;
            'd49: LUT_x2_im_res1 = 49;
            'd50: LUT_x2_im_res1 = 50;
            'd51: LUT_x2_im_res1 = 51;
            'd52: LUT_x2_im_res1 = 52;
            'd53: LUT_x2_im_res1 = 53;
            'd54: LUT_x2_im_res1 = 54;
            'd55: LUT_x2_im_res1 = 55;
            'd56: LUT_x2_im_res1 = 56;
            'd57: LUT_x2_im_res1 = 57;
            'd58: LUT_x2_im_res1 = 58;
            'd59: LUT_x2_im_res1 = 59;
            'd60: LUT_x2_im_res1 = 60;
            'd61: LUT_x2_im_res1 = 61;
            'd62: LUT_x2_im_res1 = 62;
            'd63: LUT_x2_im_res1 = 63;
            'd64: LUT_x2_im_res1 = 64;
            'd65: LUT_x2_im_res1 = 65;
            'd66: LUT_x2_im_res1 = 66;
            'd67: LUT_x2_im_res1 = 67;
            'd68: LUT_x2_im_res1 = 68;
            'd69: LUT_x2_im_res1 = 69;
            'd70: LUT_x2_im_res1 = 70;
            'd71: LUT_x2_im_res1 = 71;
            'd72: LUT_x2_im_res1 = 72;
            'd73: LUT_x2_im_res1 = 73;
            'd74: LUT_x2_im_res1 = 74;
            'd75: LUT_x2_im_res1 = 75;
            'd76: LUT_x2_im_res1 = 76;
            'd77: LUT_x2_im_res1 = 77;
            'd78: LUT_x2_im_res1 = 78;
            'd79: LUT_x2_im_res1 = 79;
            'd80: LUT_x2_im_res1 = 80;
            'd81: LUT_x2_im_res1 = 81;
            'd82: LUT_x2_im_res1 = 82;
            'd83: LUT_x2_im_res1 = 83;
            'd84: LUT_x2_im_res1 = 84;
            'd85: LUT_x2_im_res1 = 85;
            'd86: LUT_x2_im_res1 = 86;
            'd87: LUT_x2_im_res1 = 87;
            'd88: LUT_x2_im_res1 = 88;
            'd89: LUT_x2_im_res1 = 89;
            'd90: LUT_x2_im_res1 = 90;
            'd91: LUT_x2_im_res1 = 91;
            'd92: LUT_x2_im_res1 = 92;
            'd93: LUT_x2_im_res1 = 93;
            'd94: LUT_x2_im_res1 = 94;
            'd95: LUT_x2_im_res1 = 95;
            'd96: LUT_x2_im_res1 = 96;
            'd97: LUT_x2_im_res1 = 97;
            'd98: LUT_x2_im_res1 = 98;
            'd99: LUT_x2_im_res1 = 99;
            'd100: LUT_x2_im_res1 = 100;
            'd101: LUT_x2_im_res1 = 101;
            'd102: LUT_x2_im_res1 = 102;
            'd103: LUT_x2_im_res1 = 103;
            'd104: LUT_x2_im_res1 = 104;
            'd105: LUT_x2_im_res1 = 105;
            'd106: LUT_x2_im_res1 = 106;
            'd107: LUT_x2_im_res1 = 107;
            'd108: LUT_x2_im_res1 = 108;
            'd109: LUT_x2_im_res1 = 109;
            'd110: LUT_x2_im_res1 = 110;
            'd111: LUT_x2_im_res1 = 111;
            'd112: LUT_x2_im_res1 = 112;
            'd113: LUT_x2_im_res1 = 113;
            'd114: LUT_x2_im_res1 = 114;
            'd115: LUT_x2_im_res1 = 115;
            'd116: LUT_x2_im_res1 = 116;
            'd117: LUT_x2_im_res1 = 117;
            'd118: LUT_x2_im_res1 = 118;
            'd119: LUT_x2_im_res1 = 119;
            'd120: LUT_x2_im_res1 = 120;
            'd121: LUT_x2_im_res1 = 121;
            'd122: LUT_x2_im_res1 = 122;
            'd123: LUT_x2_im_res1 = 123;
            'd124: LUT_x2_im_res1 = 124;
            'd125: LUT_x2_im_res1 = 125;
            'd126: LUT_x2_im_res1 = 126;
            'd127: LUT_x2_im_res1 = 127;
            'd128: LUT_x2_im_res1 = 128;
            'd129: LUT_x2_im_res1 = 129;
            'd130: LUT_x2_im_res1 = 130;
            'd131: LUT_x2_im_res1 = 131;
            'd132: LUT_x2_im_res1 = 132;
            'd133: LUT_x2_im_res1 = 133;
            'd134: LUT_x2_im_res1 = 134;
            'd135: LUT_x2_im_res1 = 135;
            'd136: LUT_x2_im_res1 = 136;
            'd137: LUT_x2_im_res1 = 137;
            'd138: LUT_x2_im_res1 = 138;
            'd139: LUT_x2_im_res1 = 139;
            'd140: LUT_x2_im_res1 = 140;
            'd141: LUT_x2_im_res1 = 141;
            'd142: LUT_x2_im_res1 = 142;
            'd143: LUT_x2_im_res1 = 143;
            'd144: LUT_x2_im_res1 = 144;
            'd145: LUT_x2_im_res1 = 145;
            'd146: LUT_x2_im_res1 = 146;
            'd147: LUT_x2_im_res1 = 147;
            'd148: LUT_x2_im_res1 = 148;
            'd149: LUT_x2_im_res1 = 149;
            'd150: LUT_x2_im_res1 = 150;
            'd151: LUT_x2_im_res1 = 151;
            'd152: LUT_x2_im_res1 = 152;
            'd153: LUT_x2_im_res1 = 153;
            'd154: LUT_x2_im_res1 = 154;
            'd155: LUT_x2_im_res1 = 155;
            'd156: LUT_x2_im_res1 = 156;
            'd157: LUT_x2_im_res1 = 157;
            'd158: LUT_x2_im_res1 = 158;
            'd159: LUT_x2_im_res1 = 159;
            'd160: LUT_x2_im_res1 = 160;
            'd161: LUT_x2_im_res1 = 161;
            'd162: LUT_x2_im_res1 = 162;
            'd163: LUT_x2_im_res1 = 163;
            'd164: LUT_x2_im_res1 = 164;
            'd165: LUT_x2_im_res1 = 165;
            'd166: LUT_x2_im_res1 = 166;
            'd167: LUT_x2_im_res1 = 167;
            'd168: LUT_x2_im_res1 = 168;
            'd169: LUT_x2_im_res1 = 169;
            'd170: LUT_x2_im_res1 = 170;
            'd171: LUT_x2_im_res1 = 171;
            'd172: LUT_x2_im_res1 = 172;
            'd173: LUT_x2_im_res1 = 173;
            'd174: LUT_x2_im_res1 = 174;
            'd175: LUT_x2_im_res1 = 175;
            'd176: LUT_x2_im_res1 = 176;
            'd177: LUT_x2_im_res1 = 177;
            'd178: LUT_x2_im_res1 = 178;
            'd179: LUT_x2_im_res1 = 179;
            'd180: LUT_x2_im_res1 = 180;
            'd181: LUT_x2_im_res1 = 181;
            'd182: LUT_x2_im_res1 = 182;
            'd183: LUT_x2_im_res1 = 183;
            'd184: LUT_x2_im_res1 = 184;
            'd185: LUT_x2_im_res1 = 185;
            'd186: LUT_x2_im_res1 = 186;
            'd187: LUT_x2_im_res1 = 187;
            'd188: LUT_x2_im_res1 = 188;
            'd189: LUT_x2_im_res1 = 189;
            'd190: LUT_x2_im_res1 = 190;
            'd191: LUT_x2_im_res1 = 191;
            'd192: LUT_x2_im_res1 = 192;
            'd193: LUT_x2_im_res1 = 193;
            'd194: LUT_x2_im_res1 = 194;
            'd195: LUT_x2_im_res1 = 195;
            'd196: LUT_x2_im_res1 = 196;
            'd197: LUT_x2_im_res1 = 197;
            'd198: LUT_x2_im_res1 = 198;
            'd199: LUT_x2_im_res1 = 199;
            'd200: LUT_x2_im_res1 = 200;
            'd201: LUT_x2_im_res1 = 201;
            'd202: LUT_x2_im_res1 = 202;
            'd203: LUT_x2_im_res1 = 203;
            'd204: LUT_x2_im_res1 = 204;
            'd205: LUT_x2_im_res1 = 205;
            'd206: LUT_x2_im_res1 = 206;
            'd207: LUT_x2_im_res1 = 207;
            'd208: LUT_x2_im_res1 = 208;
            'd209: LUT_x2_im_res1 = 209;
            'd210: LUT_x2_im_res1 = 210;
            'd211: LUT_x2_im_res1 = 211;
            'd212: LUT_x2_im_res1 = 212;
            'd213: LUT_x2_im_res1 = 213;
            'd214: LUT_x2_im_res1 = 214;
            'd215: LUT_x2_im_res1 = 215;
            'd216: LUT_x2_im_res1 = 216;
            'd217: LUT_x2_im_res1 = 217;
            'd218: LUT_x2_im_res1 = 218;
            'd219: LUT_x2_im_res1 = 219;
            'd220: LUT_x2_im_res1 = 220;
            'd221: LUT_x2_im_res1 = 221;
            'd222: LUT_x2_im_res1 = 222;
            'd223: LUT_x2_im_res1 = 223;
            'd224: LUT_x2_im_res1 = 224;
            'd225: LUT_x2_im_res1 = 225;
            'd226: LUT_x2_im_res1 = 226;
            'd227: LUT_x2_im_res1 = 227;
            'd228: LUT_x2_im_res1 = 228;
            'd229: LUT_x2_im_res1 = 229;
            'd230: LUT_x2_im_res1 = 230;
            'd231: LUT_x2_im_res1 = 231;
            'd232: LUT_x2_im_res1 = 232;
            'd233: LUT_x2_im_res1 = 233;
            'd234: LUT_x2_im_res1 = 234;
            'd235: LUT_x2_im_res1 = 235;
            'd236: LUT_x2_im_res1 = 236;
            'd237: LUT_x2_im_res1 = 237;
            'd238: LUT_x2_im_res1 = 238;
            'd239: LUT_x2_im_res1 = 239;
            'd240: LUT_x2_im_res1 = 240;
            'd241: LUT_x2_im_res1 = 241;
            'd242: LUT_x2_im_res1 = 242;
            'd243: LUT_x2_im_res1 = 243;
            'd244: LUT_x2_im_res1 = 244;
            'd245: LUT_x2_im_res1 = 245;
            'd246: LUT_x2_im_res1 = 246;
            'd247: LUT_x2_im_res1 = 247;
            'd248: LUT_x2_im_res1 = 248;
            'd249: LUT_x2_im_res1 = 249;
            'd250: LUT_x2_im_res1 = 250;
            'd251: LUT_x2_im_res1 = 251;
            'd252: LUT_x2_im_res1 = 252;
            'd253: LUT_x2_im_res1 = 253;
            'd254: LUT_x2_im_res1 = 254;
            'd255: LUT_x2_im_res1 = 255;
            'd256: LUT_x2_im_res1 = 256;
            default: LUT_x2_im_res1 = 0;
        endcase
    end //end always */

    //X2, resonator 2, real
    always @(*) begin
        case(counter) 
            'd1: LUT_x2_real_res2 = 1;
            'd2: LUT_x2_real_res2 = 2;
            'd3: LUT_x2_real_res2 = 3;
            'd4: LUT_x2_real_res2 = 4;
            'd5: LUT_x2_real_res2 = 5;
            'd6: LUT_x2_real_res2 = 6;
            'd7: LUT_x2_real_res2 = 7;
            'd8: LUT_x2_real_res2 = 8;
            'd9: LUT_x2_real_res2 = 9;
            'd10: LUT_x2_real_res2 = 10;
            'd11: LUT_x2_real_res2 = 11;
            'd12: LUT_x2_real_res2 = 12;
            'd13: LUT_x2_real_res2 = 13;
            'd14: LUT_x2_real_res2 = 14;
            'd15: LUT_x2_real_res2 = 15;
            'd16: LUT_x2_real_res2 = 16;
            'd17: LUT_x2_real_res2 = 17;
            'd18: LUT_x2_real_res2 = 18;
            'd19: LUT_x2_real_res2 = 19;
            'd20: LUT_x2_real_res2 = 20;
            'd21: LUT_x2_real_res2 = 21;
            'd22: LUT_x2_real_res2 = 22;
            'd23: LUT_x2_real_res2 = 23;
            'd24: LUT_x2_real_res2 = 24;
            'd25: LUT_x2_real_res2 = 25;
            'd26: LUT_x2_real_res2 = 26;
            'd27: LUT_x2_real_res2 = 27;
            'd28: LUT_x2_real_res2 = 28;
            'd29: LUT_x2_real_res2 = 29;
            'd30: LUT_x2_real_res2 = 30;
            'd31: LUT_x2_real_res2 = 31;
            'd32: LUT_x2_real_res2 = 32;
            'd33: LUT_x2_real_res2 = 33;
            'd34: LUT_x2_real_res2 = 34;
            'd35: LUT_x2_real_res2 = 35;
            'd36: LUT_x2_real_res2 = 36;
            'd37: LUT_x2_real_res2 = 37;
            'd38: LUT_x2_real_res2 = 38;
            'd39: LUT_x2_real_res2 = 39;
            'd40: LUT_x2_real_res2 = 40;
            'd41: LUT_x2_real_res2 = 41;
            'd42: LUT_x2_real_res2 = 42;
            'd43: LUT_x2_real_res2 = 43;
            'd44: LUT_x2_real_res2 = 44;
            'd45: LUT_x2_real_res2 = 45;
            'd46: LUT_x2_real_res2 = 46;
            'd47: LUT_x2_real_res2 = 47;
            'd48: LUT_x2_real_res2 = 48;
            'd49: LUT_x2_real_res2 = 49;
            'd50: LUT_x2_real_res2 = 50;
            'd51: LUT_x2_real_res2 = 51;
            'd52: LUT_x2_real_res2 = 52;
            'd53: LUT_x2_real_res2 = 53;
            'd54: LUT_x2_real_res2 = 54;
            'd55: LUT_x2_real_res2 = 55;
            'd56: LUT_x2_real_res2 = 56;
            'd57: LUT_x2_real_res2 = 57;
            'd58: LUT_x2_real_res2 = 58;
            'd59: LUT_x2_real_res2 = 59;
            'd60: LUT_x2_real_res2 = 60;
            'd61: LUT_x2_real_res2 = 61;
            'd62: LUT_x2_real_res2 = 62;
            'd63: LUT_x2_real_res2 = 63;
            'd64: LUT_x2_real_res2 = 64;
            'd65: LUT_x2_real_res2 = 65;
            'd66: LUT_x2_real_res2 = 66;
            'd67: LUT_x2_real_res2 = 67;
            'd68: LUT_x2_real_res2 = 68;
            'd69: LUT_x2_real_res2 = 69;
            'd70: LUT_x2_real_res2 = 70;
            'd71: LUT_x2_real_res2 = 71;
            'd72: LUT_x2_real_res2 = 72;
            'd73: LUT_x2_real_res2 = 73;
            'd74: LUT_x2_real_res2 = 74;
            'd75: LUT_x2_real_res2 = 75;
            'd76: LUT_x2_real_res2 = 76;
            'd77: LUT_x2_real_res2 = 77;
            'd78: LUT_x2_real_res2 = 78;
            'd79: LUT_x2_real_res2 = 79;
            'd80: LUT_x2_real_res2 = 80;
            'd81: LUT_x2_real_res2 = 81;
            'd82: LUT_x2_real_res2 = 82;
            'd83: LUT_x2_real_res2 = 83;
            'd84: LUT_x2_real_res2 = 84;
            'd85: LUT_x2_real_res2 = 85;
            'd86: LUT_x2_real_res2 = 86;
            'd87: LUT_x2_real_res2 = 87;
            'd88: LUT_x2_real_res2 = 88;
            'd89: LUT_x2_real_res2 = 89;
            'd90: LUT_x2_real_res2 = 90;
            'd91: LUT_x2_real_res2 = 91;
            'd92: LUT_x2_real_res2 = 92;
            'd93: LUT_x2_real_res2 = 93;
            'd94: LUT_x2_real_res2 = 94;
            'd95: LUT_x2_real_res2 = 95;
            'd96: LUT_x2_real_res2 = 96;
            'd97: LUT_x2_real_res2 = 97;
            'd98: LUT_x2_real_res2 = 98;
            'd99: LUT_x2_real_res2 = 99;
            'd100: LUT_x2_real_res2 = 100;
            'd101: LUT_x2_real_res2 = 101;
            'd102: LUT_x2_real_res2 = 102;
            'd103: LUT_x2_real_res2 = 103;
            'd104: LUT_x2_real_res2 = 104;
            'd105: LUT_x2_real_res2 = 105;
            'd106: LUT_x2_real_res2 = 106;
            'd107: LUT_x2_real_res2 = 107;
            'd108: LUT_x2_real_res2 = 108;
            'd109: LUT_x2_real_res2 = 109;
            'd110: LUT_x2_real_res2 = 110;
            'd111: LUT_x2_real_res2 = 111;
            'd112: LUT_x2_real_res2 = 112;
            'd113: LUT_x2_real_res2 = 113;
            'd114: LUT_x2_real_res2 = 114;
            'd115: LUT_x2_real_res2 = 115;
            'd116: LUT_x2_real_res2 = 116;
            'd117: LUT_x2_real_res2 = 117;
            'd118: LUT_x2_real_res2 = 118;
            'd119: LUT_x2_real_res2 = 119;
            'd120: LUT_x2_real_res2 = 120;
            'd121: LUT_x2_real_res2 = 121;
            'd122: LUT_x2_real_res2 = 122;
            'd123: LUT_x2_real_res2 = 123;
            'd124: LUT_x2_real_res2 = 124;
            'd125: LUT_x2_real_res2 = 125;
            'd126: LUT_x2_real_res2 = 126;
            'd127: LUT_x2_real_res2 = 127;
            'd128: LUT_x2_real_res2 = 128;
            'd129: LUT_x2_real_res2 = 129;
            'd130: LUT_x2_real_res2 = 130;
            'd131: LUT_x2_real_res2 = 131;
            'd132: LUT_x2_real_res2 = 132;
            'd133: LUT_x2_real_res2 = 133;
            'd134: LUT_x2_real_res2 = 134;
            'd135: LUT_x2_real_res2 = 135;
            'd136: LUT_x2_real_res2 = 136;
            'd137: LUT_x2_real_res2 = 137;
            'd138: LUT_x2_real_res2 = 138;
            'd139: LUT_x2_real_res2 = 139;
            'd140: LUT_x2_real_res2 = 140;
            'd141: LUT_x2_real_res2 = 141;
            'd142: LUT_x2_real_res2 = 142;
            'd143: LUT_x2_real_res2 = 143;
            'd144: LUT_x2_real_res2 = 144;
            'd145: LUT_x2_real_res2 = 145;
            'd146: LUT_x2_real_res2 = 146;
            'd147: LUT_x2_real_res2 = 147;
            'd148: LUT_x2_real_res2 = 148;
            'd149: LUT_x2_real_res2 = 149;
            'd150: LUT_x2_real_res2 = 150;
            'd151: LUT_x2_real_res2 = 151;
            'd152: LUT_x2_real_res2 = 152;
            'd153: LUT_x2_real_res2 = 153;
            'd154: LUT_x2_real_res2 = 154;
            'd155: LUT_x2_real_res2 = 155;
            'd156: LUT_x2_real_res2 = 156;
            'd157: LUT_x2_real_res2 = 157;
            'd158: LUT_x2_real_res2 = 158;
            'd159: LUT_x2_real_res2 = 159;
            'd160: LUT_x2_real_res2 = 160;
            'd161: LUT_x2_real_res2 = 161;
            'd162: LUT_x2_real_res2 = 162;
            'd163: LUT_x2_real_res2 = 163;
            'd164: LUT_x2_real_res2 = 164;
            'd165: LUT_x2_real_res2 = 165;
            'd166: LUT_x2_real_res2 = 166;
            'd167: LUT_x2_real_res2 = 167;
            'd168: LUT_x2_real_res2 = 168;
            'd169: LUT_x2_real_res2 = 169;
            'd170: LUT_x2_real_res2 = 170;
            'd171: LUT_x2_real_res2 = 171;
            'd172: LUT_x2_real_res2 = 172;
            'd173: LUT_x2_real_res2 = 173;
            'd174: LUT_x2_real_res2 = 174;
            'd175: LUT_x2_real_res2 = 175;
            'd176: LUT_x2_real_res2 = 176;
            'd177: LUT_x2_real_res2 = 177;
            'd178: LUT_x2_real_res2 = 178;
            'd179: LUT_x2_real_res2 = 179;
            'd180: LUT_x2_real_res2 = 180;
            'd181: LUT_x2_real_res2 = 181;
            'd182: LUT_x2_real_res2 = 182;
            'd183: LUT_x2_real_res2 = 183;
            'd184: LUT_x2_real_res2 = 184;
            'd185: LUT_x2_real_res2 = 185;
            'd186: LUT_x2_real_res2 = 186;
            'd187: LUT_x2_real_res2 = 187;
            'd188: LUT_x2_real_res2 = 188;
            'd189: LUT_x2_real_res2 = 189;
            'd190: LUT_x2_real_res2 = 190;
            'd191: LUT_x2_real_res2 = 191;
            'd192: LUT_x2_real_res2 = 192;
            'd193: LUT_x2_real_res2 = 193;
            'd194: LUT_x2_real_res2 = 194;
            'd195: LUT_x2_real_res2 = 195;
            'd196: LUT_x2_real_res2 = 196;
            'd197: LUT_x2_real_res2 = 197;
            'd198: LUT_x2_real_res2 = 198;
            'd199: LUT_x2_real_res2 = 199;
            'd200: LUT_x2_real_res2 = 200;
            'd201: LUT_x2_real_res2 = 201;
            'd202: LUT_x2_real_res2 = 202;
            'd203: LUT_x2_real_res2 = 203;
            'd204: LUT_x2_real_res2 = 204;
            'd205: LUT_x2_real_res2 = 205;
            'd206: LUT_x2_real_res2 = 206;
            'd207: LUT_x2_real_res2 = 207;
            'd208: LUT_x2_real_res2 = 208;
            'd209: LUT_x2_real_res2 = 209;
            'd210: LUT_x2_real_res2 = 210;
            'd211: LUT_x2_real_res2 = 211;
            'd212: LUT_x2_real_res2 = 212;
            'd213: LUT_x2_real_res2 = 213;
            'd214: LUT_x2_real_res2 = 214;
            'd215: LUT_x2_real_res2 = 215;
            'd216: LUT_x2_real_res2 = 216;
            'd217: LUT_x2_real_res2 = 217;
            'd218: LUT_x2_real_res2 = 218;
            'd219: LUT_x2_real_res2 = 219;
            'd220: LUT_x2_real_res2 = 220;
            'd221: LUT_x2_real_res2 = 221;
            'd222: LUT_x2_real_res2 = 222;
            'd223: LUT_x2_real_res2 = 223;
            'd224: LUT_x2_real_res2 = 224;
            'd225: LUT_x2_real_res2 = 225;
            'd226: LUT_x2_real_res2 = 226;
            'd227: LUT_x2_real_res2 = 227;
            'd228: LUT_x2_real_res2 = 228;
            'd229: LUT_x2_real_res2 = 229;
            'd230: LUT_x2_real_res2 = 230;
            'd231: LUT_x2_real_res2 = 231;
            'd232: LUT_x2_real_res2 = 232;
            'd233: LUT_x2_real_res2 = 233;
            'd234: LUT_x2_real_res2 = 234;
            'd235: LUT_x2_real_res2 = 235;
            'd236: LUT_x2_real_res2 = 236;
            'd237: LUT_x2_real_res2 = 237;
            'd238: LUT_x2_real_res2 = 238;
            'd239: LUT_x2_real_res2 = 239;
            'd240: LUT_x2_real_res2 = 240;
            'd241: LUT_x2_real_res2 = 241;
            'd242: LUT_x2_real_res2 = 242;
            'd243: LUT_x2_real_res2 = 243;
            'd244: LUT_x2_real_res2 = 244;
            'd245: LUT_x2_real_res2 = 245;
            'd246: LUT_x2_real_res2 = 246;
            'd247: LUT_x2_real_res2 = 247;
            'd248: LUT_x2_real_res2 = 248;
            'd249: LUT_x2_real_res2 = 249;
            'd250: LUT_x2_real_res2 = 250;
            'd251: LUT_x2_real_res2 = 251;
            'd252: LUT_x2_real_res2 = 252;
            'd253: LUT_x2_real_res2 = 253;
            'd254: LUT_x2_real_res2 = 254;
            'd255: LUT_x2_real_res2 = 255;
            'd256: LUT_x2_real_res2 = 256;
            default: LUT_x2_real_res2 = 0;
        endcase
    end //end always */
    
     //X2, resonator 2, imaginary
    always @(*) begin
        case(counter) 
            'd1: LUT_x2_im_res2 = 1;
            'd2: LUT_x2_im_res2 = 2;
            'd3: LUT_x2_im_res2 = 3;
            'd4: LUT_x2_im_res2 = 4;
            'd5: LUT_x2_im_res2 = 5;
            'd6: LUT_x2_im_res2 = 6;
            'd7: LUT_x2_im_res2 = 7;
            'd8: LUT_x2_im_res2 = 8;
            'd9: LUT_x2_im_res2 = 9;
            'd10: LUT_x2_im_res2 = 10;
            'd11: LUT_x2_im_res2 = 11;
            'd12: LUT_x2_im_res2 = 12;
            'd13: LUT_x2_im_res2 = 13;
            'd14: LUT_x2_im_res2 = 14;
            'd15: LUT_x2_im_res2 = 15;
            'd16: LUT_x2_im_res2 = 16;
            'd17: LUT_x2_im_res2 = 17;
            'd18: LUT_x2_im_res2 = 18;
            'd19: LUT_x2_im_res2 = 19;
            'd20: LUT_x2_im_res2 = 20;
            'd21: LUT_x2_im_res2 = 21;
            'd22: LUT_x2_im_res2 = 22;
            'd23: LUT_x2_im_res2 = 23;
            'd24: LUT_x2_im_res2 = 24;
            'd25: LUT_x2_im_res2 = 25;
            'd26: LUT_x2_im_res2 = 26;
            'd27: LUT_x2_im_res2 = 27;
            'd28: LUT_x2_im_res2 = 28;
            'd29: LUT_x2_im_res2 = 29;
            'd30: LUT_x2_im_res2 = 30;
            'd31: LUT_x2_im_res2 = 31;
            'd32: LUT_x2_im_res2 = 32;
            'd33: LUT_x2_im_res2 = 33;
            'd34: LUT_x2_im_res2 = 34;
            'd35: LUT_x2_im_res2 = 35;
            'd36: LUT_x2_im_res2 = 36;
            'd37: LUT_x2_im_res2 = 37;
            'd38: LUT_x2_im_res2 = 38;
            'd39: LUT_x2_im_res2 = 39;
            'd40: LUT_x2_im_res2 = 40;
            'd41: LUT_x2_im_res2 = 41;
            'd42: LUT_x2_im_res2 = 42;
            'd43: LUT_x2_im_res2 = 43;
            'd44: LUT_x2_im_res2 = 44;
            'd45: LUT_x2_im_res2 = 45;
            'd46: LUT_x2_im_res2 = 46;
            'd47: LUT_x2_im_res2 = 47;
            'd48: LUT_x2_im_res2 = 48;
            'd49: LUT_x2_im_res2 = 49;
            'd50: LUT_x2_im_res2 = 50;
            'd51: LUT_x2_im_res2 = 51;
            'd52: LUT_x2_im_res2 = 52;
            'd53: LUT_x2_im_res2 = 53;
            'd54: LUT_x2_im_res2 = 54;
            'd55: LUT_x2_im_res2 = 55;
            'd56: LUT_x2_im_res2 = 56;
            'd57: LUT_x2_im_res2 = 57;
            'd58: LUT_x2_im_res2 = 58;
            'd59: LUT_x2_im_res2 = 59;
            'd60: LUT_x2_im_res2 = 60;
            'd61: LUT_x2_im_res2 = 61;
            'd62: LUT_x2_im_res2 = 62;
            'd63: LUT_x2_im_res2 = 63;
            'd64: LUT_x2_im_res2 = 64;
            'd65: LUT_x2_im_res2 = 65;
            'd66: LUT_x2_im_res2 = 66;
            'd67: LUT_x2_im_res2 = 67;
            'd68: LUT_x2_im_res2 = 68;
            'd69: LUT_x2_im_res2 = 69;
            'd70: LUT_x2_im_res2 = 70;
            'd71: LUT_x2_im_res2 = 71;
            'd72: LUT_x2_im_res2 = 72;
            'd73: LUT_x2_im_res2 = 73;
            'd74: LUT_x2_im_res2 = 74;
            'd75: LUT_x2_im_res2 = 75;
            'd76: LUT_x2_im_res2 = 76;
            'd77: LUT_x2_im_res2 = 77;
            'd78: LUT_x2_im_res2 = 78;
            'd79: LUT_x2_im_res2 = 79;
            'd80: LUT_x2_im_res2 = 80;
            'd81: LUT_x2_im_res2 = 81;
            'd82: LUT_x2_im_res2 = 82;
            'd83: LUT_x2_im_res2 = 83;
            'd84: LUT_x2_im_res2 = 84;
            'd85: LUT_x2_im_res2 = 85;
            'd86: LUT_x2_im_res2 = 86;
            'd87: LUT_x2_im_res2 = 87;
            'd88: LUT_x2_im_res2 = 88;
            'd89: LUT_x2_im_res2 = 89;
            'd90: LUT_x2_im_res2 = 90;
            'd91: LUT_x2_im_res2 = 91;
            'd92: LUT_x2_im_res2 = 92;
            'd93: LUT_x2_im_res2 = 93;
            'd94: LUT_x2_im_res2 = 94;
            'd95: LUT_x2_im_res2 = 95;
            'd96: LUT_x2_im_res2 = 96;
            'd97: LUT_x2_im_res2 = 97;
            'd98: LUT_x2_im_res2 = 98;
            'd99: LUT_x2_im_res2 = 99;
            'd100: LUT_x2_im_res2 = 100;
            'd101: LUT_x2_im_res2 = 101;
            'd102: LUT_x2_im_res2 = 102;
            'd103: LUT_x2_im_res2 = 103;
            'd104: LUT_x2_im_res2 = 104;
            'd105: LUT_x2_im_res2 = 105;
            'd106: LUT_x2_im_res2 = 106;
            'd107: LUT_x2_im_res2 = 107;
            'd108: LUT_x2_im_res2 = 108;
            'd109: LUT_x2_im_res2 = 109;
            'd110: LUT_x2_im_res2 = 110;
            'd111: LUT_x2_im_res2 = 111;
            'd112: LUT_x2_im_res2 = 112;
            'd113: LUT_x2_im_res2 = 113;
            'd114: LUT_x2_im_res2 = 114;
            'd115: LUT_x2_im_res2 = 115;
            'd116: LUT_x2_im_res2 = 116;
            'd117: LUT_x2_im_res2 = 117;
            'd118: LUT_x2_im_res2 = 118;
            'd119: LUT_x2_im_res2 = 119;
            'd120: LUT_x2_im_res2 = 120;
            'd121: LUT_x2_im_res2 = 121;
            'd122: LUT_x2_im_res2 = 122;
            'd123: LUT_x2_im_res2 = 123;
            'd124: LUT_x2_im_res2 = 124;
            'd125: LUT_x2_im_res2 = 125;
            'd126: LUT_x2_im_res2 = 126;
            'd127: LUT_x2_im_res2 = 127;
            'd128: LUT_x2_im_res2 = 128;
            'd129: LUT_x2_im_res2 = 129;
            'd130: LUT_x2_im_res2 = 130;
            'd131: LUT_x2_im_res2 = 131;
            'd132: LUT_x2_im_res2 = 132;
            'd133: LUT_x2_im_res2 = 133;
            'd134: LUT_x2_im_res2 = 134;
            'd135: LUT_x2_im_res2 = 135;
            'd136: LUT_x2_im_res2 = 136;
            'd137: LUT_x2_im_res2 = 137;
            'd138: LUT_x2_im_res2 = 138;
            'd139: LUT_x2_im_res2 = 139;
            'd140: LUT_x2_im_res2 = 140;
            'd141: LUT_x2_im_res2 = 141;
            'd142: LUT_x2_im_res2 = 142;
            'd143: LUT_x2_im_res2 = 143;
            'd144: LUT_x2_im_res2 = 144;
            'd145: LUT_x2_im_res2 = 145;
            'd146: LUT_x2_im_res2 = 146;
            'd147: LUT_x2_im_res2 = 147;
            'd148: LUT_x2_im_res2 = 148;
            'd149: LUT_x2_im_res2 = 149;
            'd150: LUT_x2_im_res2 = 150;
            'd151: LUT_x2_im_res2 = 151;
            'd152: LUT_x2_im_res2 = 152;
            'd153: LUT_x2_im_res2 = 153;
            'd154: LUT_x2_im_res2 = 154;
            'd155: LUT_x2_im_res2 = 155;
            'd156: LUT_x2_im_res2 = 156;
            'd157: LUT_x2_im_res2 = 157;
            'd158: LUT_x2_im_res2 = 158;
            'd159: LUT_x2_im_res2 = 159;
            'd160: LUT_x2_im_res2 = 160;
            'd161: LUT_x2_im_res2 = 161;
            'd162: LUT_x2_im_res2 = 162;
            'd163: LUT_x2_im_res2 = 163;
            'd164: LUT_x2_im_res2 = 164;
            'd165: LUT_x2_im_res2 = 165;
            'd166: LUT_x2_im_res2 = 166;
            'd167: LUT_x2_im_res2 = 167;
            'd168: LUT_x2_im_res2 = 168;
            'd169: LUT_x2_im_res2 = 169;
            'd170: LUT_x2_im_res2 = 170;
            'd171: LUT_x2_im_res2 = 171;
            'd172: LUT_x2_im_res2 = 172;
            'd173: LUT_x2_im_res2 = 173;
            'd174: LUT_x2_im_res2 = 174;
            'd175: LUT_x2_im_res2 = 175;
            'd176: LUT_x2_im_res2 = 176;
            'd177: LUT_x2_im_res2 = 177;
            'd178: LUT_x2_im_res2 = 178;
            'd179: LUT_x2_im_res2 = 179;
            'd180: LUT_x2_im_res2 = 180;
            'd181: LUT_x2_im_res2 = 181;
            'd182: LUT_x2_im_res2 = 182;
            'd183: LUT_x2_im_res2 = 183;
            'd184: LUT_x2_im_res2 = 184;
            'd185: LUT_x2_im_res2 = 185;
            'd186: LUT_x2_im_res2 = 186;
            'd187: LUT_x2_im_res2 = 187;
            'd188: LUT_x2_im_res2 = 188;
            'd189: LUT_x2_im_res2 = 189;
            'd190: LUT_x2_im_res2 = 190;
            'd191: LUT_x2_im_res2 = 191;
            'd192: LUT_x2_im_res2 = 192;
            'd193: LUT_x2_im_res2 = 193;
            'd194: LUT_x2_im_res2 = 194;
            'd195: LUT_x2_im_res2 = 195;
            'd196: LUT_x2_im_res2 = 196;
            'd197: LUT_x2_im_res2 = 197;
            'd198: LUT_x2_im_res2 = 198;
            'd199: LUT_x2_im_res2 = 199;
            'd200: LUT_x2_im_res2 = 200;
            'd201: LUT_x2_im_res2 = 201;
            'd202: LUT_x2_im_res2 = 202;
            'd203: LUT_x2_im_res2 = 203;
            'd204: LUT_x2_im_res2 = 204;
            'd205: LUT_x2_im_res2 = 205;
            'd206: LUT_x2_im_res2 = 206;
            'd207: LUT_x2_im_res2 = 207;
            'd208: LUT_x2_im_res2 = 208;
            'd209: LUT_x2_im_res2 = 209;
            'd210: LUT_x2_im_res2 = 210;
            'd211: LUT_x2_im_res2 = 211;
            'd212: LUT_x2_im_res2 = 212;
            'd213: LUT_x2_im_res2 = 213;
            'd214: LUT_x2_im_res2 = 214;
            'd215: LUT_x2_im_res2 = 215;
            'd216: LUT_x2_im_res2 = 216;
            'd217: LUT_x2_im_res2 = 217;
            'd218: LUT_x2_im_res2 = 218;
            'd219: LUT_x2_im_res2 = 219;
            'd220: LUT_x2_im_res2 = 220;
            'd221: LUT_x2_im_res2 = 221;
            'd222: LUT_x2_im_res2 = 222;
            'd223: LUT_x2_im_res2 = 223;
            'd224: LUT_x2_im_res2 = 224;
            'd225: LUT_x2_im_res2 = 225;
            'd226: LUT_x2_im_res2 = 226;
            'd227: LUT_x2_im_res2 = 227;
            'd228: LUT_x2_im_res2 = 228;
            'd229: LUT_x2_im_res2 = 229;
            'd230: LUT_x2_im_res2 = 230;
            'd231: LUT_x2_im_res2 = 231;
            'd232: LUT_x2_im_res2 = 232;
            'd233: LUT_x2_im_res2 = 233;
            'd234: LUT_x2_im_res2 = 234;
            'd235: LUT_x2_im_res2 = 235;
            'd236: LUT_x2_im_res2 = 236;
            'd237: LUT_x2_im_res2 = 237;
            'd238: LUT_x2_im_res2 = 238;
            'd239: LUT_x2_im_res2 = 239;
            'd240: LUT_x2_im_res2 = 240;
            'd241: LUT_x2_im_res2 = 241;
            'd242: LUT_x2_im_res2 = 242;
            'd243: LUT_x2_im_res2 = 243;
            'd244: LUT_x2_im_res2 = 244;
            'd245: LUT_x2_im_res2 = 245;
            'd246: LUT_x2_im_res2 = 246;
            'd247: LUT_x2_im_res2 = 247;
            'd248: LUT_x2_im_res2 = 248;
            'd249: LUT_x2_im_res2 = 249;
            'd250: LUT_x2_im_res2 = 250;
            'd251: LUT_x2_im_res2 = 251;
            'd252: LUT_x2_im_res2 = 252;
            'd253: LUT_x2_im_res2 = 253;
            'd254: LUT_x2_im_res2 = 254;
            'd255: LUT_x2_im_res2 = 255;
            'd256: LUT_x2_im_res2 = 256;
            default: LUT_x2_im_res2 = 0;
        endcase
    end //end always */
    
    //X3, resonator 1, real
    always @(*) begin
        case(counter) 
            'd1: LUT_x3_real_res1 = 1;
            'd2: LUT_x3_real_res1 = 2;
            'd3: LUT_x3_real_res1 = 3;
            'd4: LUT_x3_real_res1 = 4;
            'd5: LUT_x3_real_res1 = 5;
            'd6: LUT_x3_real_res1 = 6;
            'd7: LUT_x3_real_res1 = 7;
            'd8: LUT_x3_real_res1 = 8;
            'd9: LUT_x3_real_res1 = 9;
            'd10: LUT_x3_real_res1 = 10;
            'd11: LUT_x3_real_res1 = 11;
            'd12: LUT_x3_real_res1 = 12;
            'd13: LUT_x3_real_res1 = 13;
            'd14: LUT_x3_real_res1 = 14;
            'd15: LUT_x3_real_res1 = 15;
            'd16: LUT_x3_real_res1 = 16;
            'd17: LUT_x3_real_res1 = 17;
            'd18: LUT_x3_real_res1 = 18;
            'd19: LUT_x3_real_res1 = 19;
            'd20: LUT_x3_real_res1 = 20;
            'd21: LUT_x3_real_res1 = 21;
            'd22: LUT_x3_real_res1 = 22;
            'd23: LUT_x3_real_res1 = 23;
            'd24: LUT_x3_real_res1 = 24;
            'd25: LUT_x3_real_res1 = 25;
            'd26: LUT_x3_real_res1 = 26;
            'd27: LUT_x3_real_res1 = 27;
            'd28: LUT_x3_real_res1 = 28;
            'd29: LUT_x3_real_res1 = 29;
            'd30: LUT_x3_real_res1 = 30;
            'd31: LUT_x3_real_res1 = 31;
            'd32: LUT_x3_real_res1 = 32;
            'd33: LUT_x3_real_res1 = 33;
            'd34: LUT_x3_real_res1 = 34;
            'd35: LUT_x3_real_res1 = 35;
            'd36: LUT_x3_real_res1 = 36;
            'd37: LUT_x3_real_res1 = 37;
            'd38: LUT_x3_real_res1 = 38;
            'd39: LUT_x3_real_res1 = 39;
            'd40: LUT_x3_real_res1 = 40;
            'd41: LUT_x3_real_res1 = 41;
            'd42: LUT_x3_real_res1 = 42;
            'd43: LUT_x3_real_res1 = 43;
            'd44: LUT_x3_real_res1 = 44;
            'd45: LUT_x3_real_res1 = 45;
            'd46: LUT_x3_real_res1 = 46;
            'd47: LUT_x3_real_res1 = 47;
            'd48: LUT_x3_real_res1 = 48;
            'd49: LUT_x3_real_res1 = 49;
            'd50: LUT_x3_real_res1 = 50;
            'd51: LUT_x3_real_res1 = 51;
            'd52: LUT_x3_real_res1 = 52;
            'd53: LUT_x3_real_res1 = 53;
            'd54: LUT_x3_real_res1 = 54;
            'd55: LUT_x3_real_res1 = 55;
            'd56: LUT_x3_real_res1 = 56;
            'd57: LUT_x3_real_res1 = 57;
            'd58: LUT_x3_real_res1 = 58;
            'd59: LUT_x3_real_res1 = 59;
            'd60: LUT_x3_real_res1 = 60;
            'd61: LUT_x3_real_res1 = 61;
            'd62: LUT_x3_real_res1 = 62;
            'd63: LUT_x3_real_res1 = 63;
            'd64: LUT_x3_real_res1 = 64;
            'd65: LUT_x3_real_res1 = 65;
            'd66: LUT_x3_real_res1 = 66;
            'd67: LUT_x3_real_res1 = 67;
            'd68: LUT_x3_real_res1 = 68;
            'd69: LUT_x3_real_res1 = 69;
            'd70: LUT_x3_real_res1 = 70;
            'd71: LUT_x3_real_res1 = 71;
            'd72: LUT_x3_real_res1 = 72;
            'd73: LUT_x3_real_res1 = 73;
            'd74: LUT_x3_real_res1 = 74;
            'd75: LUT_x3_real_res1 = 75;
            'd76: LUT_x3_real_res1 = 76;
            'd77: LUT_x3_real_res1 = 77;
            'd78: LUT_x3_real_res1 = 78;
            'd79: LUT_x3_real_res1 = 79;
            'd80: LUT_x3_real_res1 = 80;
            'd81: LUT_x3_real_res1 = 81;
            'd82: LUT_x3_real_res1 = 82;
            'd83: LUT_x3_real_res1 = 83;
            'd84: LUT_x3_real_res1 = 84;
            'd85: LUT_x3_real_res1 = 85;
            'd86: LUT_x3_real_res1 = 86;
            'd87: LUT_x3_real_res1 = 87;
            'd88: LUT_x3_real_res1 = 88;
            'd89: LUT_x3_real_res1 = 89;
            'd90: LUT_x3_real_res1 = 90;
            'd91: LUT_x3_real_res1 = 91;
            'd92: LUT_x3_real_res1 = 92;
            'd93: LUT_x3_real_res1 = 93;
            'd94: LUT_x3_real_res1 = 94;
            'd95: LUT_x3_real_res1 = 95;
            'd96: LUT_x3_real_res1 = 96;
            'd97: LUT_x3_real_res1 = 97;
            'd98: LUT_x3_real_res1 = 98;
            'd99: LUT_x3_real_res1 = 99;
            'd100: LUT_x3_real_res1 = 100;
            'd101: LUT_x3_real_res1 = 101;
            'd102: LUT_x3_real_res1 = 102;
            'd103: LUT_x3_real_res1 = 103;
            'd104: LUT_x3_real_res1 = 104;
            'd105: LUT_x3_real_res1 = 105;
            'd106: LUT_x3_real_res1 = 106;
            'd107: LUT_x3_real_res1 = 107;
            'd108: LUT_x3_real_res1 = 108;
            'd109: LUT_x3_real_res1 = 109;
            'd110: LUT_x3_real_res1 = 110;
            'd111: LUT_x3_real_res1 = 111;
            'd112: LUT_x3_real_res1 = 112;
            'd113: LUT_x3_real_res1 = 113;
            'd114: LUT_x3_real_res1 = 114;
            'd115: LUT_x3_real_res1 = 115;
            'd116: LUT_x3_real_res1 = 116;
            'd117: LUT_x3_real_res1 = 117;
            'd118: LUT_x3_real_res1 = 118;
            'd119: LUT_x3_real_res1 = 119;
            'd120: LUT_x3_real_res1 = 120;
            'd121: LUT_x3_real_res1 = 121;
            'd122: LUT_x3_real_res1 = 122;
            'd123: LUT_x3_real_res1 = 123;
            'd124: LUT_x3_real_res1 = 124;
            'd125: LUT_x3_real_res1 = 125;
            'd126: LUT_x3_real_res1 = 126;
            'd127: LUT_x3_real_res1 = 127;
            'd128: LUT_x3_real_res1 = 128;
            'd129: LUT_x3_real_res1 = 129;
            'd130: LUT_x3_real_res1 = 130;
            'd131: LUT_x3_real_res1 = 131;
            'd132: LUT_x3_real_res1 = 132;
            'd133: LUT_x3_real_res1 = 133;
            'd134: LUT_x3_real_res1 = 134;
            'd135: LUT_x3_real_res1 = 135;
            'd136: LUT_x3_real_res1 = 136;
            'd137: LUT_x3_real_res1 = 137;
            'd138: LUT_x3_real_res1 = 138;
            'd139: LUT_x3_real_res1 = 139;
            'd140: LUT_x3_real_res1 = 140;
            'd141: LUT_x3_real_res1 = 141;
            'd142: LUT_x3_real_res1 = 142;
            'd143: LUT_x3_real_res1 = 143;
            'd144: LUT_x3_real_res1 = 144;
            'd145: LUT_x3_real_res1 = 145;
            'd146: LUT_x3_real_res1 = 146;
            'd147: LUT_x3_real_res1 = 147;
            'd148: LUT_x3_real_res1 = 148;
            'd149: LUT_x3_real_res1 = 149;
            'd150: LUT_x3_real_res1 = 150;
            'd151: LUT_x3_real_res1 = 151;
            'd152: LUT_x3_real_res1 = 152;
            'd153: LUT_x3_real_res1 = 153;
            'd154: LUT_x3_real_res1 = 154;
            'd155: LUT_x3_real_res1 = 155;
            'd156: LUT_x3_real_res1 = 156;
            'd157: LUT_x3_real_res1 = 157;
            'd158: LUT_x3_real_res1 = 158;
            'd159: LUT_x3_real_res1 = 159;
            'd160: LUT_x3_real_res1 = 160;
            'd161: LUT_x3_real_res1 = 161;
            'd162: LUT_x3_real_res1 = 162;
            'd163: LUT_x3_real_res1 = 163;
            'd164: LUT_x3_real_res1 = 164;
            'd165: LUT_x3_real_res1 = 165;
            'd166: LUT_x3_real_res1 = 166;
            'd167: LUT_x3_real_res1 = 167;
            'd168: LUT_x3_real_res1 = 168;
            'd169: LUT_x3_real_res1 = 169;
            'd170: LUT_x3_real_res1 = 170;
            'd171: LUT_x3_real_res1 = 171;
            'd172: LUT_x3_real_res1 = 172;
            'd173: LUT_x3_real_res1 = 173;
            'd174: LUT_x3_real_res1 = 174;
            'd175: LUT_x3_real_res1 = 175;
            'd176: LUT_x3_real_res1 = 176;
            'd177: LUT_x3_real_res1 = 177;
            'd178: LUT_x3_real_res1 = 178;
            'd179: LUT_x3_real_res1 = 179;
            'd180: LUT_x3_real_res1 = 180;
            'd181: LUT_x3_real_res1 = 181;
            'd182: LUT_x3_real_res1 = 182;
            'd183: LUT_x3_real_res1 = 183;
            'd184: LUT_x3_real_res1 = 184;
            'd185: LUT_x3_real_res1 = 185;
            'd186: LUT_x3_real_res1 = 186;
            'd187: LUT_x3_real_res1 = 187;
            'd188: LUT_x3_real_res1 = 188;
            'd189: LUT_x3_real_res1 = 189;
            'd190: LUT_x3_real_res1 = 190;
            'd191: LUT_x3_real_res1 = 191;
            'd192: LUT_x3_real_res1 = 192;
            'd193: LUT_x3_real_res1 = 193;
            'd194: LUT_x3_real_res1 = 194;
            'd195: LUT_x3_real_res1 = 195;
            'd196: LUT_x3_real_res1 = 196;
            'd197: LUT_x3_real_res1 = 197;
            'd198: LUT_x3_real_res1 = 198;
            'd199: LUT_x3_real_res1 = 199;
            'd200: LUT_x3_real_res1 = 200;
            'd201: LUT_x3_real_res1 = 201;
            'd202: LUT_x3_real_res1 = 202;
            'd203: LUT_x3_real_res1 = 203;
            'd204: LUT_x3_real_res1 = 204;
            'd205: LUT_x3_real_res1 = 205;
            'd206: LUT_x3_real_res1 = 206;
            'd207: LUT_x3_real_res1 = 207;
            'd208: LUT_x3_real_res1 = 208;
            'd209: LUT_x3_real_res1 = 209;
            'd210: LUT_x3_real_res1 = 210;
            'd211: LUT_x3_real_res1 = 211;
            'd212: LUT_x3_real_res1 = 212;
            'd213: LUT_x3_real_res1 = 213;
            'd214: LUT_x3_real_res1 = 214;
            'd215: LUT_x3_real_res1 = 215;
            'd216: LUT_x3_real_res1 = 216;
            'd217: LUT_x3_real_res1 = 217;
            'd218: LUT_x3_real_res1 = 218;
            'd219: LUT_x3_real_res1 = 219;
            'd220: LUT_x3_real_res1 = 220;
            'd221: LUT_x3_real_res1 = 221;
            'd222: LUT_x3_real_res1 = 222;
            'd223: LUT_x3_real_res1 = 223;
            'd224: LUT_x3_real_res1 = 224;
            'd225: LUT_x3_real_res1 = 225;
            'd226: LUT_x3_real_res1 = 226;
            'd227: LUT_x3_real_res1 = 227;
            'd228: LUT_x3_real_res1 = 228;
            'd229: LUT_x3_real_res1 = 229;
            'd230: LUT_x3_real_res1 = 230;
            'd231: LUT_x3_real_res1 = 231;
            'd232: LUT_x3_real_res1 = 232;
            'd233: LUT_x3_real_res1 = 233;
            'd234: LUT_x3_real_res1 = 234;
            'd235: LUT_x3_real_res1 = 235;
            'd236: LUT_x3_real_res1 = 236;
            'd237: LUT_x3_real_res1 = 237;
            'd238: LUT_x3_real_res1 = 238;
            'd239: LUT_x3_real_res1 = 239;
            'd240: LUT_x3_real_res1 = 240;
            'd241: LUT_x3_real_res1 = 241;
            'd242: LUT_x3_real_res1 = 242;
            'd243: LUT_x3_real_res1 = 243;
            'd244: LUT_x3_real_res1 = 244;
            'd245: LUT_x3_real_res1 = 245;
            'd246: LUT_x3_real_res1 = 246;
            'd247: LUT_x3_real_res1 = 247;
            'd248: LUT_x3_real_res1 = 248;
            'd249: LUT_x3_real_res1 = 249;
            'd250: LUT_x3_real_res1 = 250;
            'd251: LUT_x3_real_res1 = 251;
            'd252: LUT_x3_real_res1 = 252;
            'd253: LUT_x3_real_res1 = 253;
            'd254: LUT_x3_real_res1 = 254;
            'd255: LUT_x3_real_res1 = 255;
            'd256: LUT_x3_real_res1 = 256;
            default: LUT_x3_real_res1 = 0;
        endcase
    end //end always */
    
    //X3, resonator 1, imaginary
    always @(*) begin
        case(counter) 
            'd1: LUT_x3_im_res1 = 1;
            'd2: LUT_x3_im_res1 = 2;
            'd3: LUT_x3_im_res1 = 3;
            'd4: LUT_x3_im_res1 = 4;
            'd5: LUT_x3_im_res1 = 5;
            'd6: LUT_x3_im_res1 = 6;
            'd7: LUT_x3_im_res1 = 7;
            'd8: LUT_x3_im_res1 = 8;
            'd9: LUT_x3_im_res1 = 9;
            'd10: LUT_x3_im_res1 = 10;
            'd11: LUT_x3_im_res1 = 11;
            'd12: LUT_x3_im_res1 = 12;
            'd13: LUT_x3_im_res1 = 13;
            'd14: LUT_x3_im_res1 = 14;
            'd15: LUT_x3_im_res1 = 15;
            'd16: LUT_x3_im_res1 = 16;
            'd17: LUT_x3_im_res1 = 17;
            'd18: LUT_x3_im_res1 = 18;
            'd19: LUT_x3_im_res1 = 19;
            'd20: LUT_x3_im_res1 = 20;
            'd21: LUT_x3_im_res1 = 21;
            'd22: LUT_x3_im_res1 = 22;
            'd23: LUT_x3_im_res1 = 23;
            'd24: LUT_x3_im_res1 = 24;
            'd25: LUT_x3_im_res1 = 25;
            'd26: LUT_x3_im_res1 = 26;
            'd27: LUT_x3_im_res1 = 27;
            'd28: LUT_x3_im_res1 = 28;
            'd29: LUT_x3_im_res1 = 29;
            'd30: LUT_x3_im_res1 = 30;
            'd31: LUT_x3_im_res1 = 31;
            'd32: LUT_x3_im_res1 = 32;
            'd33: LUT_x3_im_res1 = 33;
            'd34: LUT_x3_im_res1 = 34;
            'd35: LUT_x3_im_res1 = 35;
            'd36: LUT_x3_im_res1 = 36;
            'd37: LUT_x3_im_res1 = 37;
            'd38: LUT_x3_im_res1 = 38;
            'd39: LUT_x3_im_res1 = 39;
            'd40: LUT_x3_im_res1 = 40;
            'd41: LUT_x3_im_res1 = 41;
            'd42: LUT_x3_im_res1 = 42;
            'd43: LUT_x3_im_res1 = 43;
            'd44: LUT_x3_im_res1 = 44;
            'd45: LUT_x3_im_res1 = 45;
            'd46: LUT_x3_im_res1 = 46;
            'd47: LUT_x3_im_res1 = 47;
            'd48: LUT_x3_im_res1 = 48;
            'd49: LUT_x3_im_res1 = 49;
            'd50: LUT_x3_im_res1 = 50;
            'd51: LUT_x3_im_res1 = 51;
            'd52: LUT_x3_im_res1 = 52;
            'd53: LUT_x3_im_res1 = 53;
            'd54: LUT_x3_im_res1 = 54;
            'd55: LUT_x3_im_res1 = 55;
            'd56: LUT_x3_im_res1 = 56;
            'd57: LUT_x3_im_res1 = 57;
            'd58: LUT_x3_im_res1 = 58;
            'd59: LUT_x3_im_res1 = 59;
            'd60: LUT_x3_im_res1 = 60;
            'd61: LUT_x3_im_res1 = 61;
            'd62: LUT_x3_im_res1 = 62;
            'd63: LUT_x3_im_res1 = 63;
            'd64: LUT_x3_im_res1 = 64;
            'd65: LUT_x3_im_res1 = 65;
            'd66: LUT_x3_im_res1 = 66;
            'd67: LUT_x3_im_res1 = 67;
            'd68: LUT_x3_im_res1 = 68;
            'd69: LUT_x3_im_res1 = 69;
            'd70: LUT_x3_im_res1 = 70;
            'd71: LUT_x3_im_res1 = 71;
            'd72: LUT_x3_im_res1 = 72;
            'd73: LUT_x3_im_res1 = 73;
            'd74: LUT_x3_im_res1 = 74;
            'd75: LUT_x3_im_res1 = 75;
            'd76: LUT_x3_im_res1 = 76;
            'd77: LUT_x3_im_res1 = 77;
            'd78: LUT_x3_im_res1 = 78;
            'd79: LUT_x3_im_res1 = 79;
            'd80: LUT_x3_im_res1 = 80;
            'd81: LUT_x3_im_res1 = 81;
            'd82: LUT_x3_im_res1 = 82;
            'd83: LUT_x3_im_res1 = 83;
            'd84: LUT_x3_im_res1 = 84;
            'd85: LUT_x3_im_res1 = 85;
            'd86: LUT_x3_im_res1 = 86;
            'd87: LUT_x3_im_res1 = 87;
            'd88: LUT_x3_im_res1 = 88;
            'd89: LUT_x3_im_res1 = 89;
            'd90: LUT_x3_im_res1 = 90;
            'd91: LUT_x3_im_res1 = 91;
            'd92: LUT_x3_im_res1 = 92;
            'd93: LUT_x3_im_res1 = 93;
            'd94: LUT_x3_im_res1 = 94;
            'd95: LUT_x3_im_res1 = 95;
            'd96: LUT_x3_im_res1 = 96;
            'd97: LUT_x3_im_res1 = 97;
            'd98: LUT_x3_im_res1 = 98;
            'd99: LUT_x3_im_res1 = 99;
            'd100: LUT_x3_im_res1 = 100;
            'd101: LUT_x3_im_res1 = 101;
            'd102: LUT_x3_im_res1 = 102;
            'd103: LUT_x3_im_res1 = 103;
            'd104: LUT_x3_im_res1 = 104;
            'd105: LUT_x3_im_res1 = 105;
            'd106: LUT_x3_im_res1 = 106;
            'd107: LUT_x3_im_res1 = 107;
            'd108: LUT_x3_im_res1 = 108;
            'd109: LUT_x3_im_res1 = 109;
            'd110: LUT_x3_im_res1 = 110;
            'd111: LUT_x3_im_res1 = 111;
            'd112: LUT_x3_im_res1 = 112;
            'd113: LUT_x3_im_res1 = 113;
            'd114: LUT_x3_im_res1 = 114;
            'd115: LUT_x3_im_res1 = 115;
            'd116: LUT_x3_im_res1 = 116;
            'd117: LUT_x3_im_res1 = 117;
            'd118: LUT_x3_im_res1 = 118;
            'd119: LUT_x3_im_res1 = 119;
            'd120: LUT_x3_im_res1 = 120;
            'd121: LUT_x3_im_res1 = 121;
            'd122: LUT_x3_im_res1 = 122;
            'd123: LUT_x3_im_res1 = 123;
            'd124: LUT_x3_im_res1 = 124;
            'd125: LUT_x3_im_res1 = 125;
            'd126: LUT_x3_im_res1 = 126;
            'd127: LUT_x3_im_res1 = 127;
            'd128: LUT_x3_im_res1 = 128;
            'd129: LUT_x3_im_res1 = 129;
            'd130: LUT_x3_im_res1 = 130;
            'd131: LUT_x3_im_res1 = 131;
            'd132: LUT_x3_im_res1 = 132;
            'd133: LUT_x3_im_res1 = 133;
            'd134: LUT_x3_im_res1 = 134;
            'd135: LUT_x3_im_res1 = 135;
            'd136: LUT_x3_im_res1 = 136;
            'd137: LUT_x3_im_res1 = 137;
            'd138: LUT_x3_im_res1 = 138;
            'd139: LUT_x3_im_res1 = 139;
            'd140: LUT_x3_im_res1 = 140;
            'd141: LUT_x3_im_res1 = 141;
            'd142: LUT_x3_im_res1 = 142;
            'd143: LUT_x3_im_res1 = 143;
            'd144: LUT_x3_im_res1 = 144;
            'd145: LUT_x3_im_res1 = 145;
            'd146: LUT_x3_im_res1 = 146;
            'd147: LUT_x3_im_res1 = 147;
            'd148: LUT_x3_im_res1 = 148;
            'd149: LUT_x3_im_res1 = 149;
            'd150: LUT_x3_im_res1 = 150;
            'd151: LUT_x3_im_res1 = 151;
            'd152: LUT_x3_im_res1 = 152;
            'd153: LUT_x3_im_res1 = 153;
            'd154: LUT_x3_im_res1 = 154;
            'd155: LUT_x3_im_res1 = 155;
            'd156: LUT_x3_im_res1 = 156;
            'd157: LUT_x3_im_res1 = 157;
            'd158: LUT_x3_im_res1 = 158;
            'd159: LUT_x3_im_res1 = 159;
            'd160: LUT_x3_im_res1 = 160;
            'd161: LUT_x3_im_res1 = 161;
            'd162: LUT_x3_im_res1 = 162;
            'd163: LUT_x3_im_res1 = 163;
            'd164: LUT_x3_im_res1 = 164;
            'd165: LUT_x3_im_res1 = 165;
            'd166: LUT_x3_im_res1 = 166;
            'd167: LUT_x3_im_res1 = 167;
            'd168: LUT_x3_im_res1 = 168;
            'd169: LUT_x3_im_res1 = 169;
            'd170: LUT_x3_im_res1 = 170;
            'd171: LUT_x3_im_res1 = 171;
            'd172: LUT_x3_im_res1 = 172;
            'd173: LUT_x3_im_res1 = 173;
            'd174: LUT_x3_im_res1 = 174;
            'd175: LUT_x3_im_res1 = 175;
            'd176: LUT_x3_im_res1 = 176;
            'd177: LUT_x3_im_res1 = 177;
            'd178: LUT_x3_im_res1 = 178;
            'd179: LUT_x3_im_res1 = 179;
            'd180: LUT_x3_im_res1 = 180;
            'd181: LUT_x3_im_res1 = 181;
            'd182: LUT_x3_im_res1 = 182;
            'd183: LUT_x3_im_res1 = 183;
            'd184: LUT_x3_im_res1 = 184;
            'd185: LUT_x3_im_res1 = 185;
            'd186: LUT_x3_im_res1 = 186;
            'd187: LUT_x3_im_res1 = 187;
            'd188: LUT_x3_im_res1 = 188;
            'd189: LUT_x3_im_res1 = 189;
            'd190: LUT_x3_im_res1 = 190;
            'd191: LUT_x3_im_res1 = 191;
            'd192: LUT_x3_im_res1 = 192;
            'd193: LUT_x3_im_res1 = 193;
            'd194: LUT_x3_im_res1 = 194;
            'd195: LUT_x3_im_res1 = 195;
            'd196: LUT_x3_im_res1 = 196;
            'd197: LUT_x3_im_res1 = 197;
            'd198: LUT_x3_im_res1 = 198;
            'd199: LUT_x3_im_res1 = 199;
            'd200: LUT_x3_im_res1 = 200;
            'd201: LUT_x3_im_res1 = 201;
            'd202: LUT_x3_im_res1 = 202;
            'd203: LUT_x3_im_res1 = 203;
            'd204: LUT_x3_im_res1 = 204;
            'd205: LUT_x3_im_res1 = 205;
            'd206: LUT_x3_im_res1 = 206;
            'd207: LUT_x3_im_res1 = 207;
            'd208: LUT_x3_im_res1 = 208;
            'd209: LUT_x3_im_res1 = 209;
            'd210: LUT_x3_im_res1 = 210;
            'd211: LUT_x3_im_res1 = 211;
            'd212: LUT_x3_im_res1 = 212;
            'd213: LUT_x3_im_res1 = 213;
            'd214: LUT_x3_im_res1 = 214;
            'd215: LUT_x3_im_res1 = 215;
            'd216: LUT_x3_im_res1 = 216;
            'd217: LUT_x3_im_res1 = 217;
            'd218: LUT_x3_im_res1 = 218;
            'd219: LUT_x3_im_res1 = 219;
            'd220: LUT_x3_im_res1 = 220;
            'd221: LUT_x3_im_res1 = 221;
            'd222: LUT_x3_im_res1 = 222;
            'd223: LUT_x3_im_res1 = 223;
            'd224: LUT_x3_im_res1 = 224;
            'd225: LUT_x3_im_res1 = 225;
            'd226: LUT_x3_im_res1 = 226;
            'd227: LUT_x3_im_res1 = 227;
            'd228: LUT_x3_im_res1 = 228;
            'd229: LUT_x3_im_res1 = 229;
            'd230: LUT_x3_im_res1 = 230;
            'd231: LUT_x3_im_res1 = 231;
            'd232: LUT_x3_im_res1 = 232;
            'd233: LUT_x3_im_res1 = 233;
            'd234: LUT_x3_im_res1 = 234;
            'd235: LUT_x3_im_res1 = 235;
            'd236: LUT_x3_im_res1 = 236;
            'd237: LUT_x3_im_res1 = 237;
            'd238: LUT_x3_im_res1 = 238;
            'd239: LUT_x3_im_res1 = 239;
            'd240: LUT_x3_im_res1 = 240;
            'd241: LUT_x3_im_res1 = 241;
            'd242: LUT_x3_im_res1 = 242;
            'd243: LUT_x3_im_res1 = 243;
            'd244: LUT_x3_im_res1 = 244;
            'd245: LUT_x3_im_res1 = 245;
            'd246: LUT_x3_im_res1 = 246;
            'd247: LUT_x3_im_res1 = 247;
            'd248: LUT_x3_im_res1 = 248;
            'd249: LUT_x3_im_res1 = 249;
            'd250: LUT_x3_im_res1 = 250;
            'd251: LUT_x3_im_res1 = 251;
            'd252: LUT_x3_im_res1 = 252;
            'd253: LUT_x3_im_res1 = 253;
            'd254: LUT_x3_im_res1 = 254;
            'd255: LUT_x3_im_res1 = 255;
            'd256: LUT_x3_im_res1 = 256;
            default: LUT_x3_im_res1 = 0;
        endcase
    end //end always */

    //X3, resonator 2, real
    always @(*) begin
        case(counter) 
            'd1: LUT_x3_real_res2 = 1;
            'd2: LUT_x3_real_res2 = 2;
            'd3: LUT_x3_real_res2 = 3;
            'd4: LUT_x3_real_res2 = 4;
            'd5: LUT_x3_real_res2 = 5;
            'd6: LUT_x3_real_res2 = 6;
            'd7: LUT_x3_real_res2 = 7;
            'd8: LUT_x3_real_res2 = 8;
            'd9: LUT_x3_real_res2 = 9;
            'd10: LUT_x3_real_res2 = 10;
            'd11: LUT_x3_real_res2 = 11;
            'd12: LUT_x3_real_res2 = 12;
            'd13: LUT_x3_real_res2 = 13;
            'd14: LUT_x3_real_res2 = 14;
            'd15: LUT_x3_real_res2 = 15;
            'd16: LUT_x3_real_res2 = 16;
            'd17: LUT_x3_real_res2 = 17;
            'd18: LUT_x3_real_res2 = 18;
            'd19: LUT_x3_real_res2 = 19;
            'd20: LUT_x3_real_res2 = 20;
            'd21: LUT_x3_real_res2 = 21;
            'd22: LUT_x3_real_res2 = 22;
            'd23: LUT_x3_real_res2 = 23;
            'd24: LUT_x3_real_res2 = 24;
            'd25: LUT_x3_real_res2 = 25;
            'd26: LUT_x3_real_res2 = 26;
            'd27: LUT_x3_real_res2 = 27;
            'd28: LUT_x3_real_res2 = 28;
            'd29: LUT_x3_real_res2 = 29;
            'd30: LUT_x3_real_res2 = 30;
            'd31: LUT_x3_real_res2 = 31;
            'd32: LUT_x3_real_res2 = 32;
            'd33: LUT_x3_real_res2 = 33;
            'd34: LUT_x3_real_res2 = 34;
            'd35: LUT_x3_real_res2 = 35;
            'd36: LUT_x3_real_res2 = 36;
            'd37: LUT_x3_real_res2 = 37;
            'd38: LUT_x3_real_res2 = 38;
            'd39: LUT_x3_real_res2 = 39;
            'd40: LUT_x3_real_res2 = 40;
            'd41: LUT_x3_real_res2 = 41;
            'd42: LUT_x3_real_res2 = 42;
            'd43: LUT_x3_real_res2 = 43;
            'd44: LUT_x3_real_res2 = 44;
            'd45: LUT_x3_real_res2 = 45;
            'd46: LUT_x3_real_res2 = 46;
            'd47: LUT_x3_real_res2 = 47;
            'd48: LUT_x3_real_res2 = 48;
            'd49: LUT_x3_real_res2 = 49;
            'd50: LUT_x3_real_res2 = 50;
            'd51: LUT_x3_real_res2 = 51;
            'd52: LUT_x3_real_res2 = 52;
            'd53: LUT_x3_real_res2 = 53;
            'd54: LUT_x3_real_res2 = 54;
            'd55: LUT_x3_real_res2 = 55;
            'd56: LUT_x3_real_res2 = 56;
            'd57: LUT_x3_real_res2 = 57;
            'd58: LUT_x3_real_res2 = 58;
            'd59: LUT_x3_real_res2 = 59;
            'd60: LUT_x3_real_res2 = 60;
            'd61: LUT_x3_real_res2 = 61;
            'd62: LUT_x3_real_res2 = 62;
            'd63: LUT_x3_real_res2 = 63;
            'd64: LUT_x3_real_res2 = 64;
            'd65: LUT_x3_real_res2 = 65;
            'd66: LUT_x3_real_res2 = 66;
            'd67: LUT_x3_real_res2 = 67;
            'd68: LUT_x3_real_res2 = 68;
            'd69: LUT_x3_real_res2 = 69;
            'd70: LUT_x3_real_res2 = 70;
            'd71: LUT_x3_real_res2 = 71;
            'd72: LUT_x3_real_res2 = 72;
            'd73: LUT_x3_real_res2 = 73;
            'd74: LUT_x3_real_res2 = 74;
            'd75: LUT_x3_real_res2 = 75;
            'd76: LUT_x3_real_res2 = 76;
            'd77: LUT_x3_real_res2 = 77;
            'd78: LUT_x3_real_res2 = 78;
            'd79: LUT_x3_real_res2 = 79;
            'd80: LUT_x3_real_res2 = 80;
            'd81: LUT_x3_real_res2 = 81;
            'd82: LUT_x3_real_res2 = 82;
            'd83: LUT_x3_real_res2 = 83;
            'd84: LUT_x3_real_res2 = 84;
            'd85: LUT_x3_real_res2 = 85;
            'd86: LUT_x3_real_res2 = 86;
            'd87: LUT_x3_real_res2 = 87;
            'd88: LUT_x3_real_res2 = 88;
            'd89: LUT_x3_real_res2 = 89;
            'd90: LUT_x3_real_res2 = 90;
            'd91: LUT_x3_real_res2 = 91;
            'd92: LUT_x3_real_res2 = 92;
            'd93: LUT_x3_real_res2 = 93;
            'd94: LUT_x3_real_res2 = 94;
            'd95: LUT_x3_real_res2 = 95;
            'd96: LUT_x3_real_res2 = 96;
            'd97: LUT_x3_real_res2 = 97;
            'd98: LUT_x3_real_res2 = 98;
            'd99: LUT_x3_real_res2 = 99;
            'd100: LUT_x3_real_res2 = 100;
            'd101: LUT_x3_real_res2 = 101;
            'd102: LUT_x3_real_res2 = 102;
            'd103: LUT_x3_real_res2 = 103;
            'd104: LUT_x3_real_res2 = 104;
            'd105: LUT_x3_real_res2 = 105;
            'd106: LUT_x3_real_res2 = 106;
            'd107: LUT_x3_real_res2 = 107;
            'd108: LUT_x3_real_res2 = 108;
            'd109: LUT_x3_real_res2 = 109;
            'd110: LUT_x3_real_res2 = 110;
            'd111: LUT_x3_real_res2 = 111;
            'd112: LUT_x3_real_res2 = 112;
            'd113: LUT_x3_real_res2 = 113;
            'd114: LUT_x3_real_res2 = 114;
            'd115: LUT_x3_real_res2 = 115;
            'd116: LUT_x3_real_res2 = 116;
            'd117: LUT_x3_real_res2 = 117;
            'd118: LUT_x3_real_res2 = 118;
            'd119: LUT_x3_real_res2 = 119;
            'd120: LUT_x3_real_res2 = 120;
            'd121: LUT_x3_real_res2 = 121;
            'd122: LUT_x3_real_res2 = 122;
            'd123: LUT_x3_real_res2 = 123;
            'd124: LUT_x3_real_res2 = 124;
            'd125: LUT_x3_real_res2 = 125;
            'd126: LUT_x3_real_res2 = 126;
            'd127: LUT_x3_real_res2 = 127;
            'd128: LUT_x3_real_res2 = 128;
            'd129: LUT_x3_real_res2 = 129;
            'd130: LUT_x3_real_res2 = 130;
            'd131: LUT_x3_real_res2 = 131;
            'd132: LUT_x3_real_res2 = 132;
            'd133: LUT_x3_real_res2 = 133;
            'd134: LUT_x3_real_res2 = 134;
            'd135: LUT_x3_real_res2 = 135;
            'd136: LUT_x3_real_res2 = 136;
            'd137: LUT_x3_real_res2 = 137;
            'd138: LUT_x3_real_res2 = 138;
            'd139: LUT_x3_real_res2 = 139;
            'd140: LUT_x3_real_res2 = 140;
            'd141: LUT_x3_real_res2 = 141;
            'd142: LUT_x3_real_res2 = 142;
            'd143: LUT_x3_real_res2 = 143;
            'd144: LUT_x3_real_res2 = 144;
            'd145: LUT_x3_real_res2 = 145;
            'd146: LUT_x3_real_res2 = 146;
            'd147: LUT_x3_real_res2 = 147;
            'd148: LUT_x3_real_res2 = 148;
            'd149: LUT_x3_real_res2 = 149;
            'd150: LUT_x3_real_res2 = 150;
            'd151: LUT_x3_real_res2 = 151;
            'd152: LUT_x3_real_res2 = 152;
            'd153: LUT_x3_real_res2 = 153;
            'd154: LUT_x3_real_res2 = 154;
            'd155: LUT_x3_real_res2 = 155;
            'd156: LUT_x3_real_res2 = 156;
            'd157: LUT_x3_real_res2 = 157;
            'd158: LUT_x3_real_res2 = 158;
            'd159: LUT_x3_real_res2 = 159;
            'd160: LUT_x3_real_res2 = 160;
            'd161: LUT_x3_real_res2 = 161;
            'd162: LUT_x3_real_res2 = 162;
            'd163: LUT_x3_real_res2 = 163;
            'd164: LUT_x3_real_res2 = 164;
            'd165: LUT_x3_real_res2 = 165;
            'd166: LUT_x3_real_res2 = 166;
            'd167: LUT_x3_real_res2 = 167;
            'd168: LUT_x3_real_res2 = 168;
            'd169: LUT_x3_real_res2 = 169;
            'd170: LUT_x3_real_res2 = 170;
            'd171: LUT_x3_real_res2 = 171;
            'd172: LUT_x3_real_res2 = 172;
            'd173: LUT_x3_real_res2 = 173;
            'd174: LUT_x3_real_res2 = 174;
            'd175: LUT_x3_real_res2 = 175;
            'd176: LUT_x3_real_res2 = 176;
            'd177: LUT_x3_real_res2 = 177;
            'd178: LUT_x3_real_res2 = 178;
            'd179: LUT_x3_real_res2 = 179;
            'd180: LUT_x3_real_res2 = 180;
            'd181: LUT_x3_real_res2 = 181;
            'd182: LUT_x3_real_res2 = 182;
            'd183: LUT_x3_real_res2 = 183;
            'd184: LUT_x3_real_res2 = 184;
            'd185: LUT_x3_real_res2 = 185;
            'd186: LUT_x3_real_res2 = 186;
            'd187: LUT_x3_real_res2 = 187;
            'd188: LUT_x3_real_res2 = 188;
            'd189: LUT_x3_real_res2 = 189;
            'd190: LUT_x3_real_res2 = 190;
            'd191: LUT_x3_real_res2 = 191;
            'd192: LUT_x3_real_res2 = 192;
            'd193: LUT_x3_real_res2 = 193;
            'd194: LUT_x3_real_res2 = 194;
            'd195: LUT_x3_real_res2 = 195;
            'd196: LUT_x3_real_res2 = 196;
            'd197: LUT_x3_real_res2 = 197;
            'd198: LUT_x3_real_res2 = 198;
            'd199: LUT_x3_real_res2 = 199;
            'd200: LUT_x3_real_res2 = 200;
            'd201: LUT_x3_real_res2 = 201;
            'd202: LUT_x3_real_res2 = 202;
            'd203: LUT_x3_real_res2 = 203;
            'd204: LUT_x3_real_res2 = 204;
            'd205: LUT_x3_real_res2 = 205;
            'd206: LUT_x3_real_res2 = 206;
            'd207: LUT_x3_real_res2 = 207;
            'd208: LUT_x3_real_res2 = 208;
            'd209: LUT_x3_real_res2 = 209;
            'd210: LUT_x3_real_res2 = 210;
            'd211: LUT_x3_real_res2 = 211;
            'd212: LUT_x3_real_res2 = 212;
            'd213: LUT_x3_real_res2 = 213;
            'd214: LUT_x3_real_res2 = 214;
            'd215: LUT_x3_real_res2 = 215;
            'd216: LUT_x3_real_res2 = 216;
            'd217: LUT_x3_real_res2 = 217;
            'd218: LUT_x3_real_res2 = 218;
            'd219: LUT_x3_real_res2 = 219;
            'd220: LUT_x3_real_res2 = 220;
            'd221: LUT_x3_real_res2 = 221;
            'd222: LUT_x3_real_res2 = 222;
            'd223: LUT_x3_real_res2 = 223;
            'd224: LUT_x3_real_res2 = 224;
            'd225: LUT_x3_real_res2 = 225;
            'd226: LUT_x3_real_res2 = 226;
            'd227: LUT_x3_real_res2 = 227;
            'd228: LUT_x3_real_res2 = 228;
            'd229: LUT_x3_real_res2 = 229;
            'd230: LUT_x3_real_res2 = 230;
            'd231: LUT_x3_real_res2 = 231;
            'd232: LUT_x3_real_res2 = 232;
            'd233: LUT_x3_real_res2 = 233;
            'd234: LUT_x3_real_res2 = 234;
            'd235: LUT_x3_real_res2 = 235;
            'd236: LUT_x3_real_res2 = 236;
            'd237: LUT_x3_real_res2 = 237;
            'd238: LUT_x3_real_res2 = 238;
            'd239: LUT_x3_real_res2 = 239;
            'd240: LUT_x3_real_res2 = 240;
            'd241: LUT_x3_real_res2 = 241;
            'd242: LUT_x3_real_res2 = 242;
            'd243: LUT_x3_real_res2 = 243;
            'd244: LUT_x3_real_res2 = 244;
            'd245: LUT_x3_real_res2 = 245;
            'd246: LUT_x3_real_res2 = 246;
            'd247: LUT_x3_real_res2 = 247;
            'd248: LUT_x3_real_res2 = 248;
            'd249: LUT_x3_real_res2 = 249;
            'd250: LUT_x3_real_res2 = 250;
            'd251: LUT_x3_real_res2 = 251;
            'd252: LUT_x3_real_res2 = 252;
            'd253: LUT_x3_real_res2 = 253;
            'd254: LUT_x3_real_res2 = 254;
            'd255: LUT_x3_real_res2 = 255;
            'd256: LUT_x3_real_res2 = 256;
            default: LUT_x3_real_res2 = 0;
        endcase
    end //end always */
    
     //X3, resonator 2, imaginary
    always @(*) begin
        case(counter) 
            'd1: LUT_x3_im_res2 = 1;
            'd2: LUT_x3_im_res2 = 2;
            'd3: LUT_x3_im_res2 = 3;
            'd4: LUT_x3_im_res2 = 4;
            'd5: LUT_x3_im_res2 = 5;
            'd6: LUT_x3_im_res2 = 6;
            'd7: LUT_x3_im_res2 = 7;
            'd8: LUT_x3_im_res2 = 8;
            'd9: LUT_x3_im_res2 = 9;
            'd10: LUT_x3_im_res2 = 10;
            'd11: LUT_x3_im_res2 = 11;
            'd12: LUT_x3_im_res2 = 12;
            'd13: LUT_x3_im_res2 = 13;
            'd14: LUT_x3_im_res2 = 14;
            'd15: LUT_x3_im_res2 = 15;
            'd16: LUT_x3_im_res2 = 16;
            'd17: LUT_x3_im_res2 = 17;
            'd18: LUT_x3_im_res2 = 18;
            'd19: LUT_x3_im_res2 = 19;
            'd20: LUT_x3_im_res2 = 20;
            'd21: LUT_x3_im_res2 = 21;
            'd22: LUT_x3_im_res2 = 22;
            'd23: LUT_x3_im_res2 = 23;
            'd24: LUT_x3_im_res2 = 24;
            'd25: LUT_x3_im_res2 = 25;
            'd26: LUT_x3_im_res2 = 26;
            'd27: LUT_x3_im_res2 = 27;
            'd28: LUT_x3_im_res2 = 28;
            'd29: LUT_x3_im_res2 = 29;
            'd30: LUT_x3_im_res2 = 30;
            'd31: LUT_x3_im_res2 = 31;
            'd32: LUT_x3_im_res2 = 32;
            'd33: LUT_x3_im_res2 = 33;
            'd34: LUT_x3_im_res2 = 34;
            'd35: LUT_x3_im_res2 = 35;
            'd36: LUT_x3_im_res2 = 36;
            'd37: LUT_x3_im_res2 = 37;
            'd38: LUT_x3_im_res2 = 38;
            'd39: LUT_x3_im_res2 = 39;
            'd40: LUT_x3_im_res2 = 40;
            'd41: LUT_x3_im_res2 = 41;
            'd42: LUT_x3_im_res2 = 42;
            'd43: LUT_x3_im_res2 = 43;
            'd44: LUT_x3_im_res2 = 44;
            'd45: LUT_x3_im_res2 = 45;
            'd46: LUT_x3_im_res2 = 46;
            'd47: LUT_x3_im_res2 = 47;
            'd48: LUT_x3_im_res2 = 48;
            'd49: LUT_x3_im_res2 = 49;
            'd50: LUT_x3_im_res2 = 50;
            'd51: LUT_x3_im_res2 = 51;
            'd52: LUT_x3_im_res2 = 52;
            'd53: LUT_x3_im_res2 = 53;
            'd54: LUT_x3_im_res2 = 54;
            'd55: LUT_x3_im_res2 = 55;
            'd56: LUT_x3_im_res2 = 56;
            'd57: LUT_x3_im_res2 = 57;
            'd58: LUT_x3_im_res2 = 58;
            'd59: LUT_x3_im_res2 = 59;
            'd60: LUT_x3_im_res2 = 60;
            'd61: LUT_x3_im_res2 = 61;
            'd62: LUT_x3_im_res2 = 62;
            'd63: LUT_x3_im_res2 = 63;
            'd64: LUT_x3_im_res2 = 64;
            'd65: LUT_x3_im_res2 = 65;
            'd66: LUT_x3_im_res2 = 66;
            'd67: LUT_x3_im_res2 = 67;
            'd68: LUT_x3_im_res2 = 68;
            'd69: LUT_x3_im_res2 = 69;
            'd70: LUT_x3_im_res2 = 70;
            'd71: LUT_x3_im_res2 = 71;
            'd72: LUT_x3_im_res2 = 72;
            'd73: LUT_x3_im_res2 = 73;
            'd74: LUT_x3_im_res2 = 74;
            'd75: LUT_x3_im_res2 = 75;
            'd76: LUT_x3_im_res2 = 76;
            'd77: LUT_x3_im_res2 = 77;
            'd78: LUT_x3_im_res2 = 78;
            'd79: LUT_x3_im_res2 = 79;
            'd80: LUT_x3_im_res2 = 80;
            'd81: LUT_x3_im_res2 = 81;
            'd82: LUT_x3_im_res2 = 82;
            'd83: LUT_x3_im_res2 = 83;
            'd84: LUT_x3_im_res2 = 84;
            'd85: LUT_x3_im_res2 = 85;
            'd86: LUT_x3_im_res2 = 86;
            'd87: LUT_x3_im_res2 = 87;
            'd88: LUT_x3_im_res2 = 88;
            'd89: LUT_x3_im_res2 = 89;
            'd90: LUT_x3_im_res2 = 90;
            'd91: LUT_x3_im_res2 = 91;
            'd92: LUT_x3_im_res2 = 92;
            'd93: LUT_x3_im_res2 = 93;
            'd94: LUT_x3_im_res2 = 94;
            'd95: LUT_x3_im_res2 = 95;
            'd96: LUT_x3_im_res2 = 96;
            'd97: LUT_x3_im_res2 = 97;
            'd98: LUT_x3_im_res2 = 98;
            'd99: LUT_x3_im_res2 = 99;
            'd100: LUT_x3_im_res2 = 100;
            'd101: LUT_x3_im_res2 = 101;
            'd102: LUT_x3_im_res2 = 102;
            'd103: LUT_x3_im_res2 = 103;
            'd104: LUT_x3_im_res2 = 104;
            'd105: LUT_x3_im_res2 = 105;
            'd106: LUT_x3_im_res2 = 106;
            'd107: LUT_x3_im_res2 = 107;
            'd108: LUT_x3_im_res2 = 108;
            'd109: LUT_x3_im_res2 = 109;
            'd110: LUT_x3_im_res2 = 110;
            'd111: LUT_x3_im_res2 = 111;
            'd112: LUT_x3_im_res2 = 112;
            'd113: LUT_x3_im_res2 = 113;
            'd114: LUT_x3_im_res2 = 114;
            'd115: LUT_x3_im_res2 = 115;
            'd116: LUT_x3_im_res2 = 116;
            'd117: LUT_x3_im_res2 = 117;
            'd118: LUT_x3_im_res2 = 118;
            'd119: LUT_x3_im_res2 = 119;
            'd120: LUT_x3_im_res2 = 120;
            'd121: LUT_x3_im_res2 = 121;
            'd122: LUT_x3_im_res2 = 122;
            'd123: LUT_x3_im_res2 = 123;
            'd124: LUT_x3_im_res2 = 124;
            'd125: LUT_x3_im_res2 = 125;
            'd126: LUT_x3_im_res2 = 126;
            'd127: LUT_x3_im_res2 = 127;
            'd128: LUT_x3_im_res2 = 128;
            'd129: LUT_x3_im_res2 = 129;
            'd130: LUT_x3_im_res2 = 130;
            'd131: LUT_x3_im_res2 = 131;
            'd132: LUT_x3_im_res2 = 132;
            'd133: LUT_x3_im_res2 = 133;
            'd134: LUT_x3_im_res2 = 134;
            'd135: LUT_x3_im_res2 = 135;
            'd136: LUT_x3_im_res2 = 136;
            'd137: LUT_x3_im_res2 = 137;
            'd138: LUT_x3_im_res2 = 138;
            'd139: LUT_x3_im_res2 = 139;
            'd140: LUT_x3_im_res2 = 140;
            'd141: LUT_x3_im_res2 = 141;
            'd142: LUT_x3_im_res2 = 142;
            'd143: LUT_x3_im_res2 = 143;
            'd144: LUT_x3_im_res2 = 144;
            'd145: LUT_x3_im_res2 = 145;
            'd146: LUT_x3_im_res2 = 146;
            'd147: LUT_x3_im_res2 = 147;
            'd148: LUT_x3_im_res2 = 148;
            'd149: LUT_x3_im_res2 = 149;
            'd150: LUT_x3_im_res2 = 150;
            'd151: LUT_x3_im_res2 = 151;
            'd152: LUT_x3_im_res2 = 152;
            'd153: LUT_x3_im_res2 = 153;
            'd154: LUT_x3_im_res2 = 154;
            'd155: LUT_x3_im_res2 = 155;
            'd156: LUT_x3_im_res2 = 156;
            'd157: LUT_x3_im_res2 = 157;
            'd158: LUT_x3_im_res2 = 158;
            'd159: LUT_x3_im_res2 = 159;
            'd160: LUT_x3_im_res2 = 160;
            'd161: LUT_x3_im_res2 = 161;
            'd162: LUT_x3_im_res2 = 162;
            'd163: LUT_x3_im_res2 = 163;
            'd164: LUT_x3_im_res2 = 164;
            'd165: LUT_x3_im_res2 = 165;
            'd166: LUT_x3_im_res2 = 166;
            'd167: LUT_x3_im_res2 = 167;
            'd168: LUT_x3_im_res2 = 168;
            'd169: LUT_x3_im_res2 = 169;
            'd170: LUT_x3_im_res2 = 170;
            'd171: LUT_x3_im_res2 = 171;
            'd172: LUT_x3_im_res2 = 172;
            'd173: LUT_x3_im_res2 = 173;
            'd174: LUT_x3_im_res2 = 174;
            'd175: LUT_x3_im_res2 = 175;
            'd176: LUT_x3_im_res2 = 176;
            'd177: LUT_x3_im_res2 = 177;
            'd178: LUT_x3_im_res2 = 178;
            'd179: LUT_x3_im_res2 = 179;
            'd180: LUT_x3_im_res2 = 180;
            'd181: LUT_x3_im_res2 = 181;
            'd182: LUT_x3_im_res2 = 182;
            'd183: LUT_x3_im_res2 = 183;
            'd184: LUT_x3_im_res2 = 184;
            'd185: LUT_x3_im_res2 = 185;
            'd186: LUT_x3_im_res2 = 186;
            'd187: LUT_x3_im_res2 = 187;
            'd188: LUT_x3_im_res2 = 188;
            'd189: LUT_x3_im_res2 = 189;
            'd190: LUT_x3_im_res2 = 190;
            'd191: LUT_x3_im_res2 = 191;
            'd192: LUT_x3_im_res2 = 192;
            'd193: LUT_x3_im_res2 = 193;
            'd194: LUT_x3_im_res2 = 194;
            'd195: LUT_x3_im_res2 = 195;
            'd196: LUT_x3_im_res2 = 196;
            'd197: LUT_x3_im_res2 = 197;
            'd198: LUT_x3_im_res2 = 198;
            'd199: LUT_x3_im_res2 = 199;
            'd200: LUT_x3_im_res2 = 200;
            'd201: LUT_x3_im_res2 = 201;
            'd202: LUT_x3_im_res2 = 202;
            'd203: LUT_x3_im_res2 = 203;
            'd204: LUT_x3_im_res2 = 204;
            'd205: LUT_x3_im_res2 = 205;
            'd206: LUT_x3_im_res2 = 206;
            'd207: LUT_x3_im_res2 = 207;
            'd208: LUT_x3_im_res2 = 208;
            'd209: LUT_x3_im_res2 = 209;
            'd210: LUT_x3_im_res2 = 210;
            'd211: LUT_x3_im_res2 = 211;
            'd212: LUT_x3_im_res2 = 212;
            'd213: LUT_x3_im_res2 = 213;
            'd214: LUT_x3_im_res2 = 214;
            'd215: LUT_x3_im_res2 = 215;
            'd216: LUT_x3_im_res2 = 216;
            'd217: LUT_x3_im_res2 = 217;
            'd218: LUT_x3_im_res2 = 218;
            'd219: LUT_x3_im_res2 = 219;
            'd220: LUT_x3_im_res2 = 220;
            'd221: LUT_x3_im_res2 = 221;
            'd222: LUT_x3_im_res2 = 222;
            'd223: LUT_x3_im_res2 = 223;
            'd224: LUT_x3_im_res2 = 224;
            'd225: LUT_x3_im_res2 = 225;
            'd226: LUT_x3_im_res2 = 226;
            'd227: LUT_x3_im_res2 = 227;
            'd228: LUT_x3_im_res2 = 228;
            'd229: LUT_x3_im_res2 = 229;
            'd230: LUT_x3_im_res2 = 230;
            'd231: LUT_x3_im_res2 = 231;
            'd232: LUT_x3_im_res2 = 232;
            'd233: LUT_x3_im_res2 = 233;
            'd234: LUT_x3_im_res2 = 234;
            'd235: LUT_x3_im_res2 = 235;
            'd236: LUT_x3_im_res2 = 236;
            'd237: LUT_x3_im_res2 = 237;
            'd238: LUT_x3_im_res2 = 238;
            'd239: LUT_x3_im_res2 = 239;
            'd240: LUT_x3_im_res2 = 240;
            'd241: LUT_x3_im_res2 = 241;
            'd242: LUT_x3_im_res2 = 242;
            'd243: LUT_x3_im_res2 = 243;
            'd244: LUT_x3_im_res2 = 244;
            'd245: LUT_x3_im_res2 = 245;
            'd246: LUT_x3_im_res2 = 246;
            'd247: LUT_x3_im_res2 = 247;
            'd248: LUT_x3_im_res2 = 248;
            'd249: LUT_x3_im_res2 = 249;
            'd250: LUT_x3_im_res2 = 250;
            'd251: LUT_x3_im_res2 = 251;
            'd252: LUT_x3_im_res2 = 252;
            'd253: LUT_x3_im_res2 = 253;
            'd254: LUT_x3_im_res2 = 254;
            'd255: LUT_x3_im_res2 = 255;
            'd256: LUT_x3_im_res2 = 256;
            default: LUT_x3_im_res2 = 0;
        endcase
    end //end always */

   
endmodule
