library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.NUMERIC_STD.ALL;

entity compare is
    generic (N : integer := 32);
    Port ( 
          
          );
end compare;

architecture behv of compare is
begin
    
end architecture;